magic
tech scmos
timestamp 1490995571
<< m2contact >>
rect -7 -7 7 7
<< end >>
