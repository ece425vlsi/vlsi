magic
tech scmos
timestamp 1493737109
<< m2contact >>
rect -2 -7 2 7
<< end >>
