magic
tech scmos
timestamp 1493747238
<< metal1 >>
rect 1178 368 1421 371
rect 346 358 909 361
rect 1106 358 1869 361
rect 178 348 869 351
rect 1050 348 1613 351
rect 30 325 2082 340
rect 55 300 2057 315
rect 55 287 2057 293
rect 540 278 550 282
rect 1082 268 1086 278
rect 450 261 461 264
rect 570 258 574 268
rect 578 258 582 267
rect 210 248 215 257
rect 226 248 230 257
rect 698 253 702 262
rect 1090 261 1094 264
rect 1109 261 1118 267
rect 1057 257 1062 261
rect 1090 258 1118 261
rect 1338 258 1342 267
rect 1418 258 1422 267
rect 818 248 823 257
rect 834 248 838 257
rect 138 234 142 242
rect 202 228 209 236
rect 250 228 254 237
rect 298 232 302 242
rect 338 228 342 237
rect 375 228 382 236
rect 418 232 422 247
rect 438 243 446 246
rect 438 241 469 243
rect 442 240 469 241
rect 503 231 510 236
rect 746 234 750 242
rect 866 238 869 253
rect 882 248 887 257
rect 930 248 934 257
rect 945 248 950 257
rect 1282 248 1286 257
rect 1010 242 1021 245
rect 1290 243 1294 252
rect 1338 250 1349 253
rect 1361 251 1374 253
rect 1361 248 1381 251
rect 1434 248 1439 257
rect 1474 248 1478 257
rect 1563 248 1573 251
rect 1594 248 1598 257
rect 1302 243 1310 246
rect 1690 243 1694 252
rect 1786 248 1790 257
rect 2002 253 2006 262
rect 1905 251 1918 253
rect 1905 248 1925 251
rect 1010 238 1014 242
rect 1302 241 1317 243
rect 1306 240 1317 241
rect 1314 231 1317 240
rect 503 228 517 231
rect 842 228 853 231
rect 1314 228 1325 231
rect 1367 228 1374 236
rect 1514 232 1518 242
rect 1554 240 1589 243
rect 1834 232 1838 242
rect 1874 228 1878 237
rect 1911 228 1915 236
rect 1021 198 1030 202
rect 1714 198 1725 201
rect 30 187 2082 193
rect 1338 178 1349 181
rect 978 158 982 168
rect 1058 158 1062 168
rect 1418 158 1422 168
rect 1682 158 1686 168
rect 474 148 485 151
rect 178 138 182 148
rect 202 138 206 148
rect 474 145 478 148
rect 783 144 790 152
rect 1114 138 1118 148
rect 1162 138 1166 147
rect 1370 144 1377 152
rect 1471 144 1478 152
rect 1730 148 1745 151
rect 1738 144 1745 148
rect 1850 141 1861 144
rect 1890 137 1901 140
rect 258 128 270 131
rect 442 130 453 133
rect 722 131 733 134
rect 1339 131 1357 134
rect 954 128 965 131
rect 1314 128 1325 131
rect 1507 128 1525 131
rect 1602 128 1606 137
rect 266 123 270 128
rect 362 125 373 128
rect 602 118 606 127
rect 650 119 655 123
rect 682 118 686 127
rect 1395 125 1405 128
rect 1274 118 1285 121
rect 1714 118 1733 121
rect 1819 119 1829 122
rect 2002 118 2006 127
rect 1714 113 1723 118
rect 1914 115 1941 118
rect 162 110 173 113
rect 493 98 509 101
rect 1202 98 1215 101
rect 55 87 2057 93
rect 55 65 2057 80
rect 30 40 2082 55
rect 42 28 757 31
rect 858 28 1453 31
rect 1458 28 1797 31
rect 602 18 1141 21
rect 1218 18 1573 21
rect 402 8 597 11
rect 914 8 1173 11
rect 1250 8 1301 11
rect 1306 8 1445 11
rect 1298 3 1301 8
rect 1466 3 1469 11
rect 1298 0 1469 3
<< metal2 >>
rect 18 377 45 380
rect 1330 379 1333 380
rect 2 268 5 321
rect 18 278 21 377
rect 1266 376 1333 379
rect 30 40 45 340
rect 55 65 70 315
rect 178 278 181 351
rect 138 238 141 271
rect 186 262 189 281
rect 186 253 190 262
rect 226 248 229 261
rect 266 243 270 252
rect 138 135 141 201
rect 170 158 173 201
rect 234 198 245 201
rect 42 0 45 31
rect 66 0 69 3
rect 98 0 101 121
rect 106 108 109 122
rect 186 118 189 134
rect 194 128 197 140
rect 202 138 205 151
rect 234 135 237 198
rect 130 108 165 111
rect 130 0 133 108
rect 170 0 173 101
rect 202 0 205 121
rect 234 0 237 131
rect 258 128 261 231
rect 266 128 269 243
rect 274 218 277 241
rect 290 178 293 264
rect 298 218 301 241
rect 306 208 309 242
rect 314 218 317 241
rect 290 138 293 151
rect 314 131 317 141
rect 266 0 269 111
rect 282 108 285 122
rect 298 109 301 131
rect 322 118 325 247
rect 330 178 333 231
rect 338 178 341 211
rect 330 138 333 151
rect 346 148 349 361
rect 354 255 357 281
rect 419 267 422 281
rect 362 247 365 261
rect 402 168 405 254
rect 434 178 437 251
rect 402 137 405 151
rect 362 108 365 128
rect 298 0 301 31
rect 330 0 333 51
rect 370 0 373 121
rect 386 98 389 117
rect 394 28 397 101
rect 410 98 413 161
rect 426 148 429 171
rect 418 118 421 141
rect 442 138 445 171
rect 450 108 453 264
rect 458 148 461 181
rect 458 78 461 101
rect 402 0 405 11
rect 434 0 437 31
rect 466 0 469 301
rect 498 281 501 361
rect 498 278 509 281
rect 546 278 549 311
rect 562 258 573 261
rect 474 98 477 242
rect 482 198 485 257
rect 586 251 589 321
rect 650 278 653 371
rect 578 248 589 251
rect 626 258 653 261
rect 490 228 493 244
rect 514 188 517 231
rect 522 191 525 231
rect 530 198 533 246
rect 546 241 557 244
rect 538 218 541 231
rect 522 188 533 191
rect 482 148 485 181
rect 490 108 493 151
rect 514 131 517 161
rect 498 0 501 61
rect 506 18 509 101
rect 522 78 525 124
rect 530 0 533 188
rect 546 181 549 241
rect 538 178 549 181
rect 554 131 557 191
rect 578 141 581 248
rect 626 247 629 258
rect 586 148 589 201
rect 602 168 605 241
rect 610 231 621 234
rect 618 181 621 231
rect 634 188 637 254
rect 642 218 645 254
rect 618 178 629 181
rect 650 178 653 258
rect 674 257 677 361
rect 658 228 661 241
rect 666 191 669 251
rect 666 188 677 191
rect 690 188 693 264
rect 730 238 733 251
rect 746 238 749 351
rect 866 331 869 351
rect 866 328 877 331
rect 778 245 781 261
rect 546 128 557 131
rect 546 8 549 128
rect 562 109 565 141
rect 578 138 589 141
rect 554 98 565 101
rect 570 98 573 131
rect 578 108 581 134
rect 586 91 589 138
rect 594 109 597 141
rect 602 138 653 141
rect 602 101 605 138
rect 570 88 589 91
rect 594 98 605 101
rect 570 0 573 88
rect 594 8 597 98
rect 618 88 621 122
rect 650 118 653 138
rect 674 115 677 188
rect 706 119 709 151
rect 722 148 725 221
rect 794 211 797 281
rect 810 235 813 311
rect 818 248 821 261
rect 826 247 829 271
rect 786 208 797 211
rect 642 81 645 112
rect 634 78 645 81
rect 602 0 605 21
rect 634 0 637 78
rect 666 0 669 101
rect 698 0 701 71
rect 730 0 733 161
rect 770 135 773 201
rect 786 148 789 208
rect 834 201 837 251
rect 858 238 869 241
rect 842 208 845 231
rect 818 198 837 201
rect 818 138 821 198
rect 810 135 821 138
rect 754 128 813 131
rect 746 109 749 121
rect 754 101 757 128
rect 738 88 741 101
rect 746 98 757 101
rect 746 78 749 98
rect 754 28 757 91
rect 762 78 765 124
rect 802 108 805 124
rect 786 88 789 101
rect 810 88 813 128
rect 826 118 829 144
rect 770 0 773 41
rect 826 38 829 101
rect 802 0 805 11
rect 834 0 837 191
rect 842 78 845 181
rect 850 158 853 201
rect 858 198 861 221
rect 866 191 869 238
rect 874 235 877 328
rect 882 248 885 271
rect 906 258 909 361
rect 890 218 893 244
rect 858 188 869 191
rect 858 126 861 188
rect 874 111 877 211
rect 882 137 885 161
rect 898 119 901 254
rect 906 228 909 241
rect 914 221 917 311
rect 1018 268 1021 311
rect 930 248 933 261
rect 906 218 917 221
rect 906 208 909 218
rect 906 198 917 201
rect 906 158 909 198
rect 858 28 861 111
rect 866 108 877 111
rect 866 0 869 108
rect 874 48 877 101
rect 898 0 901 91
rect 914 8 917 171
rect 930 127 933 161
rect 938 111 941 244
rect 946 188 949 251
rect 962 248 965 261
rect 970 248 973 264
rect 954 208 957 234
rect 994 191 997 231
rect 986 188 997 191
rect 986 148 989 188
rect 1010 181 1013 261
rect 1034 238 1037 264
rect 994 178 1013 181
rect 994 137 997 178
rect 930 108 941 111
rect 922 78 925 101
rect 930 98 933 108
rect 938 88 941 101
rect 946 78 949 122
rect 970 119 973 131
rect 1002 108 1005 141
rect 1018 118 1021 141
rect 1026 128 1029 201
rect 1042 178 1045 201
rect 1034 148 1037 161
rect 1050 151 1053 351
rect 1058 258 1061 341
rect 1066 218 1069 265
rect 1074 241 1077 291
rect 1090 198 1093 301
rect 1098 178 1101 291
rect 1106 228 1109 361
rect 1162 254 1165 311
rect 1178 278 1181 371
rect 1218 281 1221 301
rect 1186 278 1221 281
rect 1122 161 1125 254
rect 1130 208 1133 254
rect 1146 218 1149 254
rect 1210 251 1213 261
rect 1226 228 1229 241
rect 1234 221 1237 261
rect 1242 228 1245 321
rect 1266 281 1269 376
rect 1298 358 1389 361
rect 1298 328 1301 358
rect 1306 348 1381 351
rect 1306 318 1309 348
rect 1314 321 1317 341
rect 1346 321 1349 341
rect 1314 318 1349 321
rect 1250 278 1269 281
rect 1250 248 1253 278
rect 1258 251 1261 261
rect 1266 231 1269 271
rect 1258 228 1269 231
rect 1274 228 1277 291
rect 1282 248 1285 301
rect 1290 268 1293 291
rect 1226 218 1237 221
rect 1122 158 1133 161
rect 1042 148 1053 151
rect 1066 148 1101 151
rect 1034 111 1037 135
rect 1026 108 1037 111
rect 930 0 933 11
rect 970 0 973 91
rect 1018 68 1021 101
rect 1026 48 1029 108
rect 1034 41 1037 101
rect 1042 71 1045 148
rect 1050 128 1053 141
rect 1058 132 1062 142
rect 1090 108 1093 122
rect 1098 121 1101 148
rect 1114 128 1117 141
rect 1098 118 1117 121
rect 1106 101 1109 111
rect 1082 98 1109 101
rect 1042 68 1069 71
rect 1010 38 1037 41
rect 1002 0 1005 31
rect 1010 8 1013 38
rect 1034 0 1037 11
rect 1066 0 1069 68
rect 1082 38 1085 98
rect 1114 51 1117 118
rect 1122 58 1125 134
rect 1130 68 1133 158
rect 1114 48 1133 51
rect 1098 0 1101 41
rect 1130 1 1133 48
rect 1138 18 1141 171
rect 1146 118 1149 135
rect 1154 128 1157 151
rect 1210 148 1213 161
rect 1162 138 1197 141
rect 1202 128 1206 137
rect 1170 8 1173 101
rect 1178 78 1181 122
rect 1218 18 1221 201
rect 1226 168 1229 218
rect 1234 138 1237 201
rect 1258 171 1261 228
rect 1298 221 1301 252
rect 1314 241 1317 311
rect 1362 281 1365 291
rect 1322 278 1365 281
rect 1322 268 1365 271
rect 1338 258 1341 268
rect 1322 248 1341 251
rect 1354 247 1365 250
rect 1314 238 1357 241
rect 1370 231 1373 321
rect 1378 281 1381 348
rect 1386 298 1389 358
rect 1418 308 1421 371
rect 1378 278 1413 281
rect 1426 271 1429 331
rect 1410 268 1429 271
rect 1266 218 1301 221
rect 1258 168 1269 171
rect 1250 158 1261 161
rect 1250 148 1253 158
rect 1242 128 1246 137
rect 1242 81 1245 111
rect 1250 88 1253 101
rect 1258 91 1261 158
rect 1266 98 1269 168
rect 1258 88 1269 91
rect 1274 81 1277 161
rect 1282 135 1285 171
rect 1282 118 1285 131
rect 1242 78 1277 81
rect 1250 8 1253 61
rect 1282 28 1285 111
rect 1290 4 1293 141
rect 1298 81 1301 218
rect 1338 228 1373 231
rect 1338 211 1341 228
rect 1322 208 1341 211
rect 1346 208 1373 211
rect 1346 178 1349 208
rect 1306 168 1357 171
rect 1306 118 1309 168
rect 1362 161 1365 181
rect 1322 158 1365 161
rect 1314 121 1317 151
rect 1370 148 1373 208
rect 1378 168 1381 251
rect 1386 228 1389 254
rect 1410 248 1413 268
rect 1418 258 1429 261
rect 1394 239 1405 242
rect 1322 138 1365 141
rect 1322 128 1325 138
rect 1314 118 1357 121
rect 1314 111 1317 118
rect 1306 108 1317 111
rect 1330 91 1333 101
rect 1322 88 1333 91
rect 1354 88 1357 118
rect 1298 78 1309 81
rect 1306 8 1309 78
rect 1314 21 1317 71
rect 1322 61 1325 81
rect 1362 78 1365 122
rect 1386 121 1389 132
rect 1394 121 1397 239
rect 1426 235 1429 258
rect 1450 251 1453 261
rect 1434 238 1437 251
rect 1402 125 1405 211
rect 1410 138 1413 181
rect 1386 118 1397 121
rect 1322 58 1357 61
rect 1322 31 1325 51
rect 1346 31 1349 51
rect 1322 28 1349 31
rect 1362 21 1365 71
rect 1314 18 1365 21
rect 1370 8 1373 101
rect 1378 4 1381 101
rect 1418 98 1421 135
rect 1410 8 1413 91
rect 1426 88 1429 151
rect 1434 28 1437 61
rect 1442 8 1445 250
rect 1466 228 1469 246
rect 1482 231 1485 291
rect 1490 250 1493 261
rect 1498 241 1501 251
rect 1482 228 1501 231
rect 1450 28 1453 124
rect 1458 78 1461 161
rect 1474 148 1477 171
rect 1490 138 1493 161
rect 1498 125 1501 228
rect 1506 218 1509 242
rect 1514 238 1517 251
rect 1522 228 1525 264
rect 1530 251 1533 331
rect 1554 268 1557 341
rect 1538 238 1541 250
rect 1578 228 1589 231
rect 1514 148 1517 161
rect 1538 148 1541 181
rect 1578 178 1581 201
rect 1546 134 1549 161
rect 1586 158 1589 228
rect 1594 178 1597 251
rect 1602 248 1605 271
rect 1610 241 1613 351
rect 1642 257 1645 321
rect 1722 258 1757 261
rect 1602 238 1613 241
rect 1602 178 1605 238
rect 1610 208 1613 231
rect 1618 198 1621 241
rect 1458 8 1461 31
rect 1466 8 1469 91
rect 1474 38 1477 101
rect 1482 88 1485 122
rect 1554 118 1557 141
rect 1586 128 1605 131
rect 1570 18 1573 122
rect 1618 115 1621 191
rect 1626 178 1629 241
rect 1658 228 1661 241
rect 1666 228 1669 254
rect 1674 248 1693 251
rect 1674 231 1677 248
rect 1722 231 1725 258
rect 1762 251 1765 261
rect 1802 251 1805 261
rect 1674 228 1685 231
rect 1698 228 1725 231
rect 1666 151 1669 201
rect 1658 148 1669 151
rect 1650 118 1653 141
rect 1658 121 1661 148
rect 1674 118 1677 141
rect 1682 128 1685 161
rect 1690 148 1693 161
rect 1690 121 1693 135
rect 1698 128 1701 221
rect 1714 168 1717 201
rect 1698 125 1709 128
rect 1722 121 1725 228
rect 1730 208 1733 231
rect 1738 228 1741 246
rect 1746 178 1749 241
rect 1786 228 1789 251
rect 1826 228 1829 242
rect 1786 188 1789 211
rect 1730 128 1733 151
rect 1754 121 1757 132
rect 1762 123 1765 151
rect 1690 118 1725 121
rect 1730 118 1757 121
rect 1722 48 1725 101
rect 1794 28 1797 134
rect 1802 118 1805 211
rect 1842 198 1845 265
rect 1858 245 1861 301
rect 1850 181 1853 241
rect 1866 228 1869 361
rect 1890 255 1893 371
rect 1898 247 1901 361
rect 1850 178 1871 181
rect 1826 138 1829 151
rect 1826 128 1837 131
rect 1826 119 1829 128
rect 1834 118 1845 121
rect 1810 68 1813 101
rect 1834 28 1837 118
rect 1850 18 1853 144
rect 1890 137 1893 241
rect 1986 137 1989 311
rect 1986 134 1997 137
rect 1882 108 1885 124
rect 2002 118 2005 351
rect 2042 65 2057 315
rect 2067 40 2082 340
rect 1290 1 1381 4
<< metal3 >>
rect 649 367 1894 372
rect 497 357 1902 362
rect 745 347 2006 352
rect 1057 337 1318 342
rect 873 327 1302 332
rect 0 317 5 322
rect 585 317 1158 322
rect 1241 317 1310 322
rect 1153 313 1158 317
rect 1153 312 1166 313
rect 545 307 814 312
rect 913 307 1022 312
rect 1153 307 1318 312
rect 465 297 1094 302
rect 1217 297 1286 302
rect 377 287 926 292
rect 1073 287 1262 292
rect 1273 287 1294 292
rect 17 277 358 282
rect 377 277 382 287
rect 921 282 926 287
rect 1257 282 1262 287
rect 418 277 614 282
rect 793 277 918 282
rect 921 277 1182 282
rect 1257 277 1326 282
rect 913 272 918 277
rect 1 267 750 272
rect 825 267 886 272
rect 913 267 998 272
rect 1017 267 1270 272
rect 1289 267 1326 272
rect 185 257 230 262
rect 361 257 566 262
rect 577 257 702 262
rect 777 257 822 262
rect 905 257 1014 262
rect 1209 257 1262 262
rect 113 247 214 252
rect 233 247 270 252
rect 321 247 390 252
rect 409 247 438 252
rect 561 247 1110 252
rect 1137 247 1254 252
rect 1289 247 1326 252
rect 217 237 422 242
rect 521 237 662 242
rect 705 237 1078 242
rect 201 227 254 232
rect 337 227 382 232
rect 393 227 494 232
rect 521 227 1278 232
rect 273 217 646 222
rect 721 217 894 222
rect 977 217 1150 222
rect 977 212 982 217
rect 305 207 342 212
rect 401 207 846 212
rect 873 207 910 212
rect 953 207 982 212
rect 1001 207 1134 212
rect 1153 207 1326 212
rect 137 197 182 202
rect 241 197 534 202
rect 585 197 774 202
rect 849 197 982 202
rect 1001 197 1006 207
rect 1089 197 1222 202
rect 513 187 558 192
rect 633 187 822 192
rect 833 187 950 192
rect 977 182 982 197
rect 993 187 1126 192
rect 153 177 294 182
rect 310 177 334 182
rect 433 177 486 182
rect 649 177 718 182
rect 841 177 902 182
rect 977 177 1046 182
rect 249 167 406 172
rect 425 167 918 172
rect 1137 167 1230 172
rect 1281 167 1302 172
rect 169 157 710 162
rect 729 157 854 162
rect 881 157 910 162
rect 929 157 982 162
rect 1033 157 1062 162
rect 1209 157 1254 162
rect 1273 157 1326 162
rect 705 152 710 157
rect 113 147 150 152
rect 201 147 246 152
rect 289 147 334 152
rect 401 147 590 152
rect 705 147 1318 152
rect 89 137 134 142
rect 177 137 230 142
rect 273 137 598 142
rect 689 137 854 142
rect 897 137 1326 142
rect 129 132 134 137
rect 129 127 198 132
rect 233 127 302 132
rect 337 127 446 132
rect 481 127 574 132
rect 609 127 958 132
rect 969 127 1054 132
rect 1113 127 1158 132
rect 1201 127 1286 132
rect 81 117 102 122
rect 185 117 326 122
rect 369 117 686 122
rect 745 117 1022 122
rect 1145 117 1294 122
rect 1305 112 1310 122
rect 105 107 134 112
rect 209 107 286 112
rect 361 107 494 112
rect 537 107 1094 112
rect 1105 107 1246 112
rect 1281 107 1310 112
rect 361 102 366 107
rect 1321 102 1326 112
rect 169 97 366 102
rect 385 97 414 102
rect 473 97 934 102
rect 1017 97 1206 102
rect 1265 97 1326 102
rect 65 87 742 92
rect 753 87 790 92
rect 809 87 862 92
rect 897 87 942 92
rect 969 87 1254 92
rect 1265 87 1326 92
rect 65 0 70 87
rect 857 82 862 87
rect 457 77 526 82
rect 641 77 750 82
rect 761 77 846 82
rect 857 77 926 82
rect 945 77 1030 82
rect 1177 77 1326 82
rect 697 67 1022 72
rect 1129 67 1318 72
rect 497 57 1254 62
rect 329 47 878 52
rect 1025 47 1326 52
rect 769 37 830 42
rect 849 37 1086 42
rect 1097 37 1326 42
rect 1330 40 1336 340
rect 1345 337 1558 342
rect 1425 327 1534 332
rect 1369 317 1646 322
rect 1339 65 1345 315
rect 1417 307 1990 312
rect 1385 297 1862 302
rect 1361 287 1486 292
rect 1361 267 1454 272
rect 1529 267 1606 272
rect 1449 262 1454 267
rect 1393 257 1422 262
rect 1449 257 1806 262
rect 1361 247 1414 252
rect 1441 247 1478 252
rect 1497 247 1518 252
rect 1569 247 1710 252
rect 1921 247 1998 252
rect 1353 237 1390 242
rect 1433 237 1542 242
rect 1617 237 1686 242
rect 1745 237 1782 242
rect 1809 237 1838 242
rect 1865 237 1894 242
rect 1385 232 1390 237
rect 1385 227 1582 232
rect 1625 227 1670 232
rect 1681 227 1830 232
rect 1873 227 1915 232
rect 1441 217 1702 222
rect 1401 207 1478 212
rect 1593 207 1734 212
rect 1801 207 1942 212
rect 1577 197 1622 202
rect 1649 197 1846 202
rect 1617 187 1790 192
rect 1361 177 1630 182
rect 1353 167 1382 172
rect 1473 167 1718 172
rect 1417 157 1462 162
rect 1489 157 1550 162
rect 1585 157 1694 162
rect 1665 147 1766 152
rect 1785 147 1905 152
rect 1361 137 1830 142
rect 1521 127 1590 132
rect 1641 127 1734 132
rect 1833 127 1878 132
rect 1393 117 1542 122
rect 1553 117 1678 122
rect 1801 117 1846 122
rect 1449 107 1942 112
rect 1377 97 1638 102
rect 1721 97 1788 102
rect 1353 87 1414 92
rect 1425 87 1486 92
rect 1361 77 1462 82
rect 1361 67 1814 72
rect 1353 57 1438 62
rect 1345 47 1726 52
rect 849 32 854 37
rect 1321 32 1326 37
rect 1345 37 1478 42
rect 1345 32 1350 37
rect 297 27 398 32
rect 433 27 854 32
rect 1001 27 1286 32
rect 1321 27 1350 32
rect 1433 27 1838 32
rect 505 17 1854 22
rect 545 7 806 12
rect 929 7 1014 12
rect 1033 7 1374 12
rect 1409 7 1462 12
use $$M3_M2  $$M3_M2_0
timestamp 1493737109
transform 1 0 652 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1493737109
transform 1 0 1180 0 1 370
box -2 -2 2 2
use $$M2_M1  $$M2_M1_1
timestamp 1493737109
transform 1 0 1420 0 1 370
box -2 -2 2 2
use $$M3_M2  $$M3_M2_1
timestamp 1493737109
transform 1 0 1892 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1493737109
transform 1 0 348 0 1 360
box -2 -2 2 2
use $$M3_M2  $$M3_M2_2
timestamp 1493737109
transform 1 0 500 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_3
timestamp 1493737109
transform 1 0 676 0 1 360
box -2 -2 2 2
use $$M2_M1  $$M2_M1_4
timestamp 1493737109
transform 1 0 908 0 1 360
box -2 -2 2 2
use $$M2_M1  $$M2_M1_5
timestamp 1493737109
transform 1 0 1108 0 1 360
box -2 -2 2 2
use $$M2_M1  $$M2_M1_6
timestamp 1493737109
transform 1 0 1868 0 1 360
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1493737109
transform 1 0 1900 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_7
timestamp 1493737109
transform 1 0 180 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1493737109
transform 1 0 748 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_8
timestamp 1493737109
transform 1 0 868 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_9
timestamp 1493737109
transform 1 0 1052 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_10
timestamp 1493737109
transform 1 0 1612 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_5
timestamp 1493737109
transform 1 0 2004 0 1 350
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1493737109
transform 1 0 37 0 1 332
box -7 -7 7 7
use $$M3_M2  $$M3_M2_6
timestamp 1493737109
transform 1 0 1060 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_7
timestamp 1493737109
transform 1 0 1316 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_8
timestamp 1493737109
transform 1 0 1348 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_9
timestamp 1493737109
transform 1 0 1556 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_10
timestamp 1493737109
transform 1 0 876 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_11
timestamp 1493737109
transform 1 0 1300 0 1 330
box -3 -3 3 3
use $$M3_M2_1500_1500_1_2  $$M3_M2_1500_1500_1_2_0
timestamp 1493737109
transform 1 0 1333 0 1 332
box -3 -6 3 5
use $$M3_M2  $$M3_M2_12
timestamp 1493737109
transform 1 0 1428 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_13
timestamp 1493737109
transform 1 0 1532 0 1 330
box -3 -3 3 3
use $$M2_M1_1500_1500_1_3  $$M2_M1_1500_1500_1_3_0
timestamp 1493737109
transform 1 0 1333 0 1 332
box -2 -7 2 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1493737109
transform 1 0 2074 0 1 332
box -7 -7 7 7
use $$M3_M2  $$M3_M2_14
timestamp 1493737109
transform 1 0 4 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_15
timestamp 1493737109
transform 1 0 588 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_16
timestamp 1493737109
transform 1 0 1244 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_17
timestamp 1493737109
transform 1 0 1308 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_18
timestamp 1493737109
transform 1 0 1372 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_19
timestamp 1493737109
transform 1 0 1644 0 1 320
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1493737109
transform 1 0 62 0 1 307
box -7 -7 7 7
use $$M3_M2  $$M3_M2_20
timestamp 1493737109
transform 1 0 548 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1493737109
transform 1 0 812 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_22
timestamp 1493737109
transform 1 0 916 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_23
timestamp 1493737109
transform 1 0 1020 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_24
timestamp 1493737109
transform 1 0 1164 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_25
timestamp 1493737109
transform 1 0 1316 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_28
timestamp 1493737109
transform 1 0 468 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_29
timestamp 1493737109
transform 1 0 1092 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_30
timestamp 1493737109
transform 1 0 1220 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_31
timestamp 1493737109
transform 1 0 1284 0 1 300
box -3 -3 3 3
use $$M3_M2_1500_1500_1_2  $$M3_M2_1500_1500_1_2_1
timestamp 1493737109
transform 1 0 1342 0 1 307
box -3 -6 3 5
use $$M3_M2  $$M3_M2_26
timestamp 1493737109
transform 1 0 1420 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_27
timestamp 1493737109
transform 1 0 1988 0 1 310
box -3 -3 3 3
use $$M2_M1_1500_1500_1_3  $$M2_M1_1500_1500_1_3_1
timestamp 1493737109
transform 1 0 1342 0 1 307
box -2 -7 2 7
use $$M3_M2  $$M3_M2_32
timestamp 1493737109
transform 1 0 1388 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_33
timestamp 1493737109
transform 1 0 1860 0 1 300
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1493737109
transform 1 0 2049 0 1 307
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1493737109
transform 1 0 62 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_34
timestamp 1493737109
transform 1 0 20 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1493737109
transform 1 0 180 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_36
timestamp 1493737109
transform 1 0 4 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_37
timestamp 1493737109
transform 1 0 140 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_38
timestamp 1493737109
transform 1 0 116 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_12
timestamp 1493737109
transform 1 0 116 0 1 246
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1493737109
transform 1 0 140 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_35
timestamp 1493737109
transform 1 0 188 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_39
timestamp 1493737109
transform 1 0 188 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_14
timestamp 1493737109
transform 1 0 188 0 1 255
box -2 -2 2 2
use $$M3_M2  $$M3_M2_40
timestamp 1493737109
transform 1 0 140 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_15
timestamp 1493737109
transform 1 0 172 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_16
timestamp 1493737109
transform 1 0 180 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_41
timestamp 1493737109
transform 1 0 180 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_42
timestamp 1493737109
transform 1 0 228 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_18
timestamp 1493737109
transform 1 0 212 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_43
timestamp 1493737109
transform 1 0 212 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_19
timestamp 1493737109
transform 1 0 228 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_17
timestamp 1493737109
transform 1 0 236 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1493737109
transform 1 0 236 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_20
timestamp 1493737109
transform 1 0 220 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_45
timestamp 1493737109
transform 1 0 220 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_21
timestamp 1493737109
transform 1 0 204 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_46
timestamp 1493737109
transform 1 0 204 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_47
timestamp 1493737109
transform 1 0 268 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_22
timestamp 1493737109
transform 1 0 268 0 1 245
box -2 -2 2 2
use $$M2_M1  $$M2_M1_24
timestamp 1493737109
transform 1 0 252 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1493737109
transform 1 0 252 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_23
timestamp 1493737109
transform 1 0 276 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_25
timestamp 1493737109
transform 1 0 260 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_26
timestamp 1493737109
transform 1 0 244 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_50
timestamp 1493737109
transform 1 0 244 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_49
timestamp 1493737109
transform 1 0 276 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_27
timestamp 1493737109
transform 1 0 292 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_51
timestamp 1493737109
transform 1 0 324 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_28
timestamp 1493737109
transform 1 0 324 0 1 246
box -2 -2 2 2
use $$M2_M1  $$M2_M1_30
timestamp 1493737109
transform 1 0 300 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_29
timestamp 1493737109
transform 1 0 308 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_31
timestamp 1493737109
transform 1 0 316 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_32
timestamp 1493737109
transform 1 0 332 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_53
timestamp 1493737109
transform 1 0 300 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_54
timestamp 1493737109
transform 1 0 316 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_55
timestamp 1493737109
transform 1 0 308 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_33
timestamp 1493737109
transform 1 0 340 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_52
timestamp 1493737109
transform 1 0 340 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_56
timestamp 1493737109
transform 1 0 340 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_57
timestamp 1493737109
transform 1 0 356 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_34
timestamp 1493737109
transform 1 0 380 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_58
timestamp 1493737109
transform 1 0 380 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_35
timestamp 1493737109
transform 1 0 356 0 1 257
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1493737109
transform 1 0 364 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_36
timestamp 1493737109
transform 1 0 364 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_37
timestamp 1493737109
transform 1 0 388 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_38
timestamp 1493737109
transform 1 0 404 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_64
timestamp 1493737109
transform 1 0 421 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_41
timestamp 1493737109
transform 1 0 421 0 1 269
box -2 -2 2 2
use $$M3_M2  $$M3_M2_60
timestamp 1493737109
transform 1 0 388 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_39
timestamp 1493737109
transform 1 0 380 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_61
timestamp 1493737109
transform 1 0 380 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_43
timestamp 1493737109
transform 1 0 412 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_65
timestamp 1493737109
transform 1 0 412 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1493737109
transform 1 0 436 0 1 251
box -2 -2 2 2
use $$M3_M2  $$M3_M2_66
timestamp 1493737109
transform 1 0 436 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_40
timestamp 1493737109
transform 1 0 396 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1493737109
transform 1 0 396 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_63
timestamp 1493737109
transform 1 0 404 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_45
timestamp 1493737109
transform 1 0 420 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_67
timestamp 1493737109
transform 1 0 420 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_42
timestamp 1493737109
transform 1 0 452 0 1 263
box -2 -2 2 2
use $$M2_M1  $$M2_M1_47
timestamp 1493737109
transform 1 0 484 0 1 256
box -2 -2 2 2
use $$M2_M1  $$M2_M1_46
timestamp 1493737109
transform 1 0 508 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1493737109
transform 1 0 476 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_48
timestamp 1493737109
transform 1 0 492 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_68
timestamp 1493737109
transform 1 0 492 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_69
timestamp 1493737109
transform 1 0 484 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_50
timestamp 1493737109
transform 1 0 548 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_51
timestamp 1493737109
transform 1 0 532 0 1 245
box -2 -2 2 2
use $$M3_M2  $$M3_M2_70
timestamp 1493737109
transform 1 0 564 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_52
timestamp 1493737109
transform 1 0 572 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_53
timestamp 1493737109
transform 1 0 580 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_71
timestamp 1493737109
transform 1 0 580 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1493737109
transform 1 0 564 0 1 251
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1493737109
transform 1 0 564 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_56
timestamp 1493737109
transform 1 0 524 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_73
timestamp 1493737109
transform 1 0 524 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_57
timestamp 1493737109
transform 1 0 516 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_74
timestamp 1493737109
transform 1 0 524 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_55
timestamp 1493737109
transform 1 0 556 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_58
timestamp 1493737109
transform 1 0 540 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_75
timestamp 1493737109
transform 1 0 540 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_76
timestamp 1493737109
transform 1 0 532 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_60
timestamp 1493737109
transform 1 0 588 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_79
timestamp 1493737109
transform 1 0 588 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1493737109
transform 1 0 596 0 1 259
box -2 -2 2 2
use $$M3_M2  $$M3_M2_77
timestamp 1493737109
transform 1 0 596 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1493737109
transform 1 0 612 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_80
timestamp 1493737109
transform 1 0 612 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_78
timestamp 1493737109
transform 1 0 604 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_62
timestamp 1493737109
transform 1 0 652 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_63
timestamp 1493737109
transform 1 0 636 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_64
timestamp 1493737109
transform 1 0 644 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_65
timestamp 1493737109
transform 1 0 628 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_66
timestamp 1493737109
transform 1 0 612 0 1 233
box -2 -2 2 2
use $$M2_M1  $$M2_M1_67
timestamp 1493737109
transform 1 0 676 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_68
timestamp 1493737109
transform 1 0 668 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_81
timestamp 1493737109
transform 1 0 660 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_69
timestamp 1493737109
transform 1 0 660 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_82
timestamp 1493737109
transform 1 0 644 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_70
timestamp 1493737109
transform 1 0 692 0 1 263
box -2 -2 2 2
use $$M2_M1  $$M2_M1_71
timestamp 1493737109
transform 1 0 700 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_83
timestamp 1493737109
transform 1 0 700 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_84
timestamp 1493737109
transform 1 0 796 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_85
timestamp 1493737109
transform 1 0 748 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_86
timestamp 1493737109
transform 1 0 780 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_87
timestamp 1493737109
transform 1 0 732 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_72
timestamp 1493737109
transform 1 0 780 0 1 247
box -2 -2 2 2
use $$M2_M1  $$M2_M1_73
timestamp 1493737109
transform 1 0 708 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_88
timestamp 1493737109
transform 1 0 708 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_74
timestamp 1493737109
transform 1 0 732 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_75
timestamp 1493737109
transform 1 0 748 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_89
timestamp 1493737109
transform 1 0 828 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_90
timestamp 1493737109
transform 1 0 820 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_76
timestamp 1493737109
transform 1 0 820 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_78
timestamp 1493737109
transform 1 0 828 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_77
timestamp 1493737109
transform 1 0 836 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_79
timestamp 1493737109
transform 1 0 812 0 1 237
box -2 -2 2 2
use $$M3_M2  $$M3_M2_91
timestamp 1493737109
transform 1 0 724 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_92
timestamp 1493737109
transform 1 0 772 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_81
timestamp 1493737109
transform 1 0 844 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_97
timestamp 1493737109
transform 1 0 844 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_93
timestamp 1493737109
transform 1 0 860 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_80
timestamp 1493737109
transform 1 0 868 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_94
timestamp 1493737109
transform 1 0 884 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_95
timestamp 1493737109
transform 1 0 908 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_83
timestamp 1493737109
transform 1 0 884 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_82
timestamp 1493737109
transform 1 0 900 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_84
timestamp 1493737109
transform 1 0 892 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_85
timestamp 1493737109
transform 1 0 876 0 1 237
box -2 -2 2 2
use $$M3_M2  $$M3_M2_96
timestamp 1493737109
transform 1 0 860 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_101
timestamp 1493737109
transform 1 0 852 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_98
timestamp 1493737109
transform 1 0 908 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_86
timestamp 1493737109
transform 1 0 908 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_99
timestamp 1493737109
transform 1 0 892 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_100
timestamp 1493737109
transform 1 0 876 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_87
timestamp 1493737109
transform 1 0 860 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_102
timestamp 1493737109
transform 1 0 908 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_103
timestamp 1493737109
transform 1 0 932 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_88
timestamp 1493737109
transform 1 0 924 0 1 251
box -2 -2 2 2
use $$M3_M2  $$M3_M2_105
timestamp 1493737109
transform 1 0 964 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_93
timestamp 1493737109
transform 1 0 972 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_104
timestamp 1493737109
transform 1 0 924 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_89
timestamp 1493737109
transform 1 0 932 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_90
timestamp 1493737109
transform 1 0 948 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_91
timestamp 1493737109
transform 1 0 916 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_92
timestamp 1493737109
transform 1 0 940 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_94
timestamp 1493737109
transform 1 0 964 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_95
timestamp 1493737109
transform 1 0 956 0 1 233
box -2 -2 2 2
use $$M3_M2  $$M3_M2_107
timestamp 1493737109
transform 1 0 956 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_106
timestamp 1493737109
transform 1 0 972 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_96
timestamp 1493737109
transform 1 0 996 0 1 270
box -2 -2 2 2
use $$M3_M2  $$M3_M2_108
timestamp 1493737109
transform 1 0 996 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_109
timestamp 1493737109
transform 1 0 1020 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_110
timestamp 1493737109
transform 1 0 1012 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_97
timestamp 1493737109
transform 1 0 1004 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_111
timestamp 1493737109
transform 1 0 1004 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_98
timestamp 1493737109
transform 1 0 1012 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_99
timestamp 1493737109
transform 1 0 996 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_100
timestamp 1493737109
transform 1 0 1004 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_112
timestamp 1493737109
transform 1 0 1004 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_101
timestamp 1493737109
transform 1 0 1036 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_113
timestamp 1493737109
transform 1 0 1076 0 1 290
box -3 -3 3 3
use $$M2_M1  $$M2_M1_102
timestamp 1493737109
transform 1 0 1084 0 1 270
box -2 -2 2 2
use $$M3_M2  $$M3_M2_115
timestamp 1493737109
transform 1 0 1084 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_103
timestamp 1493737109
transform 1 0 1068 0 1 264
box -2 -2 2 2
use $$M2_M1  $$M2_M1_104
timestamp 1493737109
transform 1 0 1060 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_116
timestamp 1493737109
transform 1 0 1036 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_105
timestamp 1493737109
transform 1 0 1028 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_106
timestamp 1493737109
transform 1 0 1044 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_107
timestamp 1493737109
transform 1 0 1076 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_117
timestamp 1493737109
transform 1 0 1076 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_118
timestamp 1493737109
transform 1 0 1068 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_114
timestamp 1493737109
transform 1 0 1100 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_119
timestamp 1493737109
transform 1 0 1092 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_120
timestamp 1493737109
transform 1 0 1108 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_110
timestamp 1493737109
transform 1 0 1108 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_108
timestamp 1493737109
transform 1 0 1124 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_109
timestamp 1493737109
transform 1 0 1132 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_111
timestamp 1493737109
transform 1 0 1116 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_121
timestamp 1493737109
transform 1 0 1116 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_122
timestamp 1493737109
transform 1 0 1132 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_113
timestamp 1493737109
transform 1 0 1140 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_112
timestamp 1493737109
transform 1 0 1148 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_123
timestamp 1493737109
transform 1 0 1140 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_124
timestamp 1493737109
transform 1 0 1148 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_125
timestamp 1493737109
transform 1 0 1180 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_114
timestamp 1493737109
transform 1 0 1188 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_115
timestamp 1493737109
transform 1 0 1164 0 1 256
box -2 -2 2 2
use $$M2_M1  $$M2_M1_117
timestamp 1493737109
transform 1 0 1156 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_127
timestamp 1493737109
transform 1 0 1156 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_126
timestamp 1493737109
transform 1 0 1212 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_116
timestamp 1493737109
transform 1 0 1212 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_133
timestamp 1493737109
transform 1 0 1276 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_134
timestamp 1493737109
transform 1 0 1292 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_135
timestamp 1493737109
transform 1 0 1268 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_136
timestamp 1493737109
transform 1 0 1292 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_128
timestamp 1493737109
transform 1 0 1236 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_129
timestamp 1493737109
transform 1 0 1260 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_130
timestamp 1493737109
transform 1 0 1252 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_118
timestamp 1493737109
transform 1 0 1260 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_119
timestamp 1493737109
transform 1 0 1236 0 1 245
box -2 -2 2 2
use $$M2_M1  $$M2_M1_120
timestamp 1493737109
transform 1 0 1228 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_131
timestamp 1493737109
transform 1 0 1228 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_121
timestamp 1493737109
transform 1 0 1244 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_132
timestamp 1493737109
transform 1 0 1220 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_122
timestamp 1493737109
transform 1 0 1236 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_124
timestamp 1493737109
transform 1 0 1284 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_125
timestamp 1493737109
transform 1 0 1292 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_123
timestamp 1493737109
transform 1 0 1300 0 1 251
box -2 -2 2 2
use $$M3_M2  $$M3_M2_137
timestamp 1493737109
transform 1 0 1292 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_126
timestamp 1493737109
transform 1 0 1276 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_138
timestamp 1493737109
transform 1 0 1276 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_127
timestamp 1493737109
transform 1 0 1268 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_141
timestamp 1493737109
transform 1 0 1324 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_142
timestamp 1493737109
transform 1 0 1324 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_144
timestamp 1493737109
transform 1 0 1324 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_131
timestamp 1493737109
transform 1 0 1324 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_146
timestamp 1493737109
transform 1 0 1324 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_128
timestamp 1493737109
transform 1 0 1342 0 1 290
box -2 -2 2 2
use $$M3_M2  $$M3_M2_139
timestamp 1493737109
transform 1 0 1342 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_140
timestamp 1493737109
transform 1 0 1364 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_143
timestamp 1493737109
transform 1 0 1364 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_129
timestamp 1493737109
transform 1 0 1340 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_130
timestamp 1493737109
transform 1 0 1340 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_132
timestamp 1493737109
transform 1 0 1356 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_145
timestamp 1493737109
transform 1 0 1364 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_147
timestamp 1493737109
transform 1 0 1356 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_133
timestamp 1493737109
transform 1 0 1372 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_134
timestamp 1493737109
transform 1 0 1412 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_135
timestamp 1493737109
transform 1 0 1396 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_148
timestamp 1493737109
transform 1 0 1396 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_136
timestamp 1493737109
transform 1 0 1420 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_149
timestamp 1493737109
transform 1 0 1420 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_138
timestamp 1493737109
transform 1 0 1380 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_137
timestamp 1493737109
transform 1 0 1388 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_150
timestamp 1493737109
transform 1 0 1412 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_139
timestamp 1493737109
transform 1 0 1404 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_151
timestamp 1493737109
transform 1 0 1388 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_152
timestamp 1493737109
transform 1 0 1404 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_153
timestamp 1493737109
transform 1 0 1452 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_141
timestamp 1493737109
transform 1 0 1436 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_142
timestamp 1493737109
transform 1 0 1444 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_154
timestamp 1493737109
transform 1 0 1444 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_140
timestamp 1493737109
transform 1 0 1452 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_143
timestamp 1493737109
transform 1 0 1428 0 1 237
box -2 -2 2 2
use $$M3_M2  $$M3_M2_155
timestamp 1493737109
transform 1 0 1436 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_156
timestamp 1493737109
transform 1 0 1444 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_157
timestamp 1493737109
transform 1 0 1484 0 1 290
box -3 -3 3 3
use $$M3_M2  $$M3_M2_158
timestamp 1493737109
transform 1 0 1492 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_148
timestamp 1493737109
transform 1 0 1476 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_144
timestamp 1493737109
transform 1 0 1492 0 1 252
box -2 -2 2 2
use $$M3_M2  $$M3_M2_159
timestamp 1493737109
transform 1 0 1532 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_145
timestamp 1493737109
transform 1 0 1556 0 1 270
box -2 -2 2 2
use $$M2_M1  $$M2_M1_146
timestamp 1493737109
transform 1 0 1524 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_160
timestamp 1493737109
transform 1 0 1476 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_161
timestamp 1493737109
transform 1 0 1500 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_162
timestamp 1493737109
transform 1 0 1516 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_147
timestamp 1493737109
transform 1 0 1532 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_149
timestamp 1493737109
transform 1 0 1468 0 1 244
box -2 -2 2 2
use $$M3_M2  $$M3_M2_163
timestamp 1493737109
transform 1 0 1468 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_150
timestamp 1493737109
transform 1 0 1500 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_151
timestamp 1493737109
transform 1 0 1508 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_152
timestamp 1493737109
transform 1 0 1516 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_164
timestamp 1493737109
transform 1 0 1508 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_153
timestamp 1493737109
transform 1 0 1476 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_165
timestamp 1493737109
transform 1 0 1476 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_155
timestamp 1493737109
transform 1 0 1540 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_167
timestamp 1493737109
transform 1 0 1540 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_168
timestamp 1493737109
transform 1 0 1524 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_154
timestamp 1493737109
transform 1 0 1572 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_166
timestamp 1493737109
transform 1 0 1572 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_158
timestamp 1493737109
transform 1 0 1580 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_170
timestamp 1493737109
transform 1 0 1580 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_175
timestamp 1493737109
transform 1 0 1580 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_169
timestamp 1493737109
transform 1 0 1604 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_156
timestamp 1493737109
transform 1 0 1596 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_157
timestamp 1493737109
transform 1 0 1604 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_159
timestamp 1493737109
transform 1 0 1620 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_171
timestamp 1493737109
transform 1 0 1620 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_160
timestamp 1493737109
transform 1 0 1628 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_161
timestamp 1493737109
transform 1 0 1612 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_172
timestamp 1493737109
transform 1 0 1628 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_173
timestamp 1493737109
transform 1 0 1596 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_174
timestamp 1493737109
transform 1 0 1612 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_176
timestamp 1493737109
transform 1 0 1620 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_162
timestamp 1493737109
transform 1 0 1644 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_163
timestamp 1493737109
transform 1 0 1668 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_164
timestamp 1493737109
transform 1 0 1676 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_165
timestamp 1493737109
transform 1 0 1692 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_178
timestamp 1493737109
transform 1 0 1660 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_167
timestamp 1493737109
transform 1 0 1684 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_179
timestamp 1493737109
transform 1 0 1684 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_168
timestamp 1493737109
transform 1 0 1660 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_180
timestamp 1493737109
transform 1 0 1668 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_181
timestamp 1493737109
transform 1 0 1684 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_166
timestamp 1493737109
transform 1 0 1708 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_177
timestamp 1493737109
transform 1 0 1708 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_169
timestamp 1493737109
transform 1 0 1700 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_170
timestamp 1493737109
transform 1 0 1652 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_182
timestamp 1493737109
transform 1 0 1652 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_183
timestamp 1493737109
transform 1 0 1668 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_184
timestamp 1493737109
transform 1 0 1700 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_176
timestamp 1493737109
transform 1 0 1716 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_171
timestamp 1493737109
transform 1 0 1756 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_172
timestamp 1493737109
transform 1 0 1740 0 1 245
box -2 -2 2 2
use $$M3_M2  $$M3_M2_185
timestamp 1493737109
transform 1 0 1764 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_173
timestamp 1493737109
transform 1 0 1764 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_174
timestamp 1493737109
transform 1 0 1748 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_186
timestamp 1493737109
transform 1 0 1748 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_175
timestamp 1493737109
transform 1 0 1732 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_187
timestamp 1493737109
transform 1 0 1740 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_188
timestamp 1493737109
transform 1 0 1732 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_189
timestamp 1493737109
transform 1 0 1804 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_178
timestamp 1493737109
transform 1 0 1788 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_177
timestamp 1493737109
transform 1 0 1804 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_180
timestamp 1493737109
transform 1 0 1780 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_190
timestamp 1493737109
transform 1 0 1780 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_179
timestamp 1493737109
transform 1 0 1812 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_191
timestamp 1493737109
transform 1 0 1812 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_192
timestamp 1493737109
transform 1 0 1788 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_181
timestamp 1493737109
transform 1 0 1788 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_193
timestamp 1493737109
transform 1 0 1804 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_182
timestamp 1493737109
transform 1 0 1844 0 1 264
box -2 -2 2 2
use $$M2_M1  $$M2_M1_183
timestamp 1493737109
transform 1 0 1828 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_185
timestamp 1493737109
transform 1 0 1836 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_194
timestamp 1493737109
transform 1 0 1836 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_184
timestamp 1493737109
transform 1 0 1860 0 1 247
box -2 -2 2 2
use $$M2_M1  $$M2_M1_186
timestamp 1493737109
transform 1 0 1852 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_196
timestamp 1493737109
transform 1 0 1828 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_195
timestamp 1493737109
transform 1 0 1868 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_187
timestamp 1493737109
transform 1 0 1868 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_198
timestamp 1493737109
transform 1 0 1844 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_188
timestamp 1493737109
transform 1 0 1876 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_197
timestamp 1493737109
transform 1 0 1876 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_189
timestamp 1493737109
transform 1 0 1892 0 1 257
box -2 -2 2 2
use $$M2_M1  $$M2_M1_192
timestamp 1493737109
transform 1 0 1900 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_201
timestamp 1493737109
transform 1 0 1892 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_191
timestamp 1493737109
transform 1 0 1924 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_199
timestamp 1493737109
transform 1 0 1924 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_193
timestamp 1493737109
transform 1 0 1913 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_202
timestamp 1493737109
transform 1 0 1913 0 1 230
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1493737109
transform 1 0 2049 0 1 290
box -7 -2 7 2
use $$M2_M1  $$M2_M1_190
timestamp 1493737109
transform 1 0 2004 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_200
timestamp 1493737109
transform 1 0 1996 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_194
timestamp 1493737109
transform 1 0 1996 0 1 246
box -2 -2 2 2
use $$M2_M1  $$M2_M1_195
timestamp 1493737109
transform 1 0 1940 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_203
timestamp 1493737109
transform 1 0 1940 0 1 210
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1493737109
transform 1 0 37 0 1 190
box -7 -2 7 2
use DFFPOSX1  DFFPOSX1_0
timestamp 1493737109
transform 1 0 80 0 -1 290
box -8 -3 104 105
use INVX2  INVX2_0
timestamp 1493737109
transform -1 0 192 0 -1 290
box -9 -3 26 105
use FILL  FILL_0
timestamp 1493737109
transform 1 0 192 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1493737109
transform -1 0 232 0 -1 290
box -8 -3 34 105
use INVX2  INVX2_1
timestamp 1493737109
transform 1 0 232 0 -1 290
box -9 -3 26 105
use NAND3X1  NAND3X1_0
timestamp 1493737109
transform -1 0 280 0 -1 290
box -8 -3 40 105
use FILL  FILL_1
timestamp 1493737109
transform 1 0 280 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1493737109
transform 1 0 288 0 -1 290
box -8 -3 32 105
use NAND3X1  NAND3X1_1
timestamp 1493737109
transform 1 0 312 0 -1 290
box -8 -3 40 105
use FILL  FILL_2
timestamp 1493737109
transform 1 0 344 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1493737109
transform 1 0 352 0 -1 290
box -8 -3 34 105
use INVX2  INVX2_2
timestamp 1493737109
transform 1 0 384 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1493737109
transform 1 0 400 0 -1 290
box -9 -3 26 105
use AOI21X1  AOI21X1_0
timestamp 1493737109
transform -1 0 448 0 -1 290
box -7 -3 39 105
use FILL  FILL_3
timestamp 1493737109
transform 1 0 448 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1493737109
transform 1 0 456 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_204
timestamp 1493737109
transform 1 0 516 0 1 190
box -3 -3 3 3
use OAI21X1  OAI21X1_2
timestamp 1493737109
transform 1 0 480 0 -1 290
box -8 -3 34 105
use FILL  FILL_4
timestamp 1493737109
transform 1 0 512 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_205
timestamp 1493737109
transform 1 0 556 0 1 190
box -3 -3 3 3
use NAND3X1  NAND3X1_2
timestamp 1493737109
transform 1 0 520 0 -1 290
box -8 -3 40 105
use AOI21X1  AOI21X1_1
timestamp 1493737109
transform 1 0 552 0 -1 290
box -7 -3 39 105
use INVX2  INVX2_4
timestamp 1493737109
transform -1 0 600 0 -1 290
box -9 -3 26 105
use FILL  FILL_5
timestamp 1493737109
transform 1 0 600 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_206
timestamp 1493737109
transform 1 0 636 0 1 190
box -3 -3 3 3
use OAI21X1  OAI21X1_3
timestamp 1493737109
transform -1 0 640 0 -1 290
box -8 -3 34 105
use $$M3_M2  $$M3_M2_207
timestamp 1493737109
transform 1 0 668 0 1 190
box -3 -3 3 3
use INVX2  INVX2_5
timestamp 1493737109
transform 1 0 640 0 -1 290
box -9 -3 26 105
use NAND2X1  NAND2X1_0
timestamp 1493737109
transform -1 0 680 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_208
timestamp 1493737109
transform 1 0 692 0 1 190
box -3 -3 3 3
use FILL  FILL_6
timestamp 1493737109
transform 1 0 680 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1493737109
transform 1 0 688 0 -1 290
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_1
timestamp 1493737109
transform -1 0 808 0 -1 290
box -8 -3 104 105
use $$M3_M2  $$M3_M2_209
timestamp 1493737109
transform 1 0 820 0 1 190
box -3 -3 3 3
use $$M3_M2  $$M3_M2_210
timestamp 1493737109
transform 1 0 836 0 1 190
box -3 -3 3 3
use OAI21X1  OAI21X1_4
timestamp 1493737109
transform -1 0 840 0 -1 290
box -8 -3 34 105
use FILL  FILL_7
timestamp 1493737109
transform 1 0 840 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1493737109
transform -1 0 872 0 -1 290
box -8 -3 32 105
use OAI21X1  OAI21X1_5
timestamp 1493737109
transform -1 0 904 0 -1 290
box -8 -3 34 105
use NAND2X1  NAND2X1_2
timestamp 1493737109
transform -1 0 928 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_211
timestamp 1493737109
transform 1 0 948 0 1 190
box -3 -3 3 3
use OAI21X1  OAI21X1_6
timestamp 1493737109
transform 1 0 928 0 -1 290
box -8 -3 34 105
use INVX1  INVX1_0
timestamp 1493737109
transform -1 0 976 0 -1 290
box -9 -3 26 105
use FILL  FILL_8
timestamp 1493737109
transform 1 0 976 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_212
timestamp 1493737109
transform 1 0 996 0 1 190
box -3 -3 3 3
use NAND3X1  NAND3X1_3
timestamp 1493737109
transform -1 0 1016 0 -1 290
box -8 -3 40 105
use NOR2X1  NOR2X1_3
timestamp 1493737109
transform -1 0 1040 0 -1 290
box -8 -3 32 105
use OR2X1  OR2X1_0
timestamp 1493737109
transform -1 0 1072 0 -1 290
box -8 -3 40 105
use NOR2X1  NOR2X1_4
timestamp 1493737109
transform -1 0 1096 0 -1 290
box -8 -3 32 105
use FILL  FILL_9
timestamp 1493737109
transform 1 0 1096 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_213
timestamp 1493737109
transform 1 0 1124 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_3
timestamp 1493737109
transform -1 0 1128 0 -1 290
box -8 -3 32 105
use INVX2  INVX2_6
timestamp 1493737109
transform 1 0 1128 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1493737109
transform 1 0 1144 0 -1 290
box -9 -3 26 105
use XOR2X1  XOR2X1_0
timestamp 1493737109
transform 1 0 1160 0 -1 290
box -8 -3 64 105
use FILL  FILL_10
timestamp 1493737109
transform 1 0 1216 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1493737109
transform 1 0 1224 0 -1 290
box -8 -3 40 105
use INVX2  INVX2_8
timestamp 1493737109
transform 1 0 1256 0 -1 290
box -9 -3 26 105
use AOI22X1  AOI22X1_0
timestamp 1493737109
transform -1 0 1312 0 -1 290
box -8 -3 46 105
use FILL  FILL_11
timestamp 1493737109
transform 1 0 1312 0 -1 290
box -8 -3 16 105
use $$M2_M1  $$M2_M1_196
timestamp 1493737109
transform 1 0 1333 0 1 190
box -2 -2 2 2
use $$M3_M2  $$M3_M2_214
timestamp 1493737109
transform 1 0 1333 0 1 190
box -3 -3 3 3
use NOR2X1  NOR2X1_5
timestamp 1493737109
transform -1 0 1344 0 -1 290
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1493737109
transform 1 0 1344 0 -1 290
box -8 -3 34 105
use FILL  FILL_12
timestamp 1493737109
transform 1 0 1376 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1493737109
transform 1 0 1384 0 -1 290
box -9 -3 26 105
use NOR2X1  NOR2X1_6
timestamp 1493737109
transform -1 0 1424 0 -1 290
box -8 -3 32 105
use OAI21X1  OAI21X1_8
timestamp 1493737109
transform -1 0 1456 0 -1 290
box -8 -3 34 105
use FILL  FILL_13
timestamp 1493737109
transform 1 0 1456 0 -1 290
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1493737109
transform -1 0 1504 0 -1 290
box -8 -3 46 105
use NOR2X1  NOR2X1_7
timestamp 1493737109
transform -1 0 1528 0 -1 290
box -8 -3 32 105
use OAI22X1  OAI22X1_0
timestamp 1493737109
transform 1 0 1528 0 -1 290
box -8 -3 46 105
use FILL  FILL_14
timestamp 1493737109
transform 1 0 1568 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1493737109
transform -1 0 1600 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_215
timestamp 1493737109
transform 1 0 1620 0 1 190
box -3 -3 3 3
use NAND3X1  NAND3X1_5
timestamp 1493737109
transform -1 0 1632 0 -1 290
box -8 -3 40 105
use FILL  FILL_15
timestamp 1493737109
transform 1 0 1632 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1493737109
transform 1 0 1640 0 -1 290
box -8 -3 32 105
use INVX2  INVX2_10
timestamp 1493737109
transform 1 0 1664 0 -1 290
box -9 -3 26 105
use NAND3X1  NAND3X1_6
timestamp 1493737109
transform 1 0 1680 0 -1 290
box -8 -3 40 105
use FILL  FILL_16
timestamp 1493737109
transform 1 0 1712 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1493737109
transform -1 0 1752 0 -1 290
box -8 -3 40 105
use INVX2  INVX2_11
timestamp 1493737109
transform -1 0 1768 0 -1 290
box -9 -3 26 105
use FILL  FILL_17
timestamp 1493737109
transform 1 0 1768 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_216
timestamp 1493737109
transform 1 0 1788 0 1 190
box -3 -3 3 3
use AOI22X1  AOI22X1_2
timestamp 1493737109
transform -1 0 1816 0 -1 290
box -8 -3 46 105
use FILL  FILL_18
timestamp 1493737109
transform 1 0 1816 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1493737109
transform -1 0 1848 0 -1 290
box -8 -3 32 105
use NAND3X1  NAND3X1_8
timestamp 1493737109
transform 1 0 1848 0 -1 290
box -8 -3 40 105
use FILL  FILL_19
timestamp 1493737109
transform 1 0 1880 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1493737109
transform 1 0 1888 0 -1 290
box -8 -3 34 105
use FILL  FILL_20
timestamp 1493737109
transform 1 0 1920 0 -1 290
box -8 -3 16 105
use FILL  FILL_21
timestamp 1493737109
transform 1 0 1928 0 -1 290
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_2
timestamp 1493737109
transform -1 0 2032 0 -1 290
box -8 -3 104 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1493737109
transform 1 0 2074 0 1 190
box -7 -2 7 2
use $$M2_M1  $$M2_M1_197
timestamp 1493737109
transform 1 0 92 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_217
timestamp 1493737109
transform 1 0 92 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_198
timestamp 1493737109
transform 1 0 84 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_218
timestamp 1493737109
transform 1 0 84 0 1 120
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1493737109
transform 1 0 62 0 1 90
box -7 -2 7 2
use $$M2_M1  $$M2_M1_199
timestamp 1493737109
transform 1 0 116 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_219
timestamp 1493737109
transform 1 0 116 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_220
timestamp 1493737109
transform 1 0 100 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_200
timestamp 1493737109
transform 1 0 108 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_221
timestamp 1493737109
transform 1 0 108 0 1 110
box -3 -3 3 3
use INVX2  INVX2_12
timestamp 1493737109
transform 1 0 80 0 1 90
box -9 -3 26 105
use FILL  FILL_22
timestamp 1493737109
transform -1 0 104 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_201
timestamp 1493737109
transform 1 0 156 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_222
timestamp 1493737109
transform 1 0 156 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_202
timestamp 1493737109
transform 1 0 148 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_223
timestamp 1493737109
transform 1 0 148 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_203
timestamp 1493737109
transform 1 0 132 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_224
timestamp 1493737109
transform 1 0 132 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_204
timestamp 1493737109
transform 1 0 140 0 1 137
box -2 -2 2 2
use $$M3_M2  $$M3_M2_228
timestamp 1493737109
transform 1 0 132 0 1 110
box -3 -3 3 3
use INVX2  INVX2_13
timestamp 1493737109
transform 1 0 104 0 1 90
box -9 -3 26 105
use FILL  FILL_23
timestamp 1493737109
transform -1 0 128 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_225
timestamp 1493737109
transform 1 0 172 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_207
timestamp 1493737109
transform 1 0 164 0 1 110
box -2 -2 2 2
use NAND3X1  NAND3X1_9
timestamp 1493737109
transform 1 0 128 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_205
timestamp 1493737109
transform 1 0 180 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_226
timestamp 1493737109
transform 1 0 180 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_227
timestamp 1493737109
transform 1 0 204 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_208
timestamp 1493737109
transform 1 0 196 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_206
timestamp 1493737109
transform 1 0 204 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_232
timestamp 1493737109
transform 1 0 172 0 1 100
box -3 -3 3 3
use FILL  FILL_24
timestamp 1493737109
transform -1 0 168 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_209
timestamp 1493737109
transform 1 0 188 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_229
timestamp 1493737109
transform 1 0 196 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_230
timestamp 1493737109
transform 1 0 188 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_231
timestamp 1493737109
transform 1 0 204 0 1 120
box -3 -3 3 3
use NOR2X1  NOR2X1_9
timestamp 1493737109
transform 1 0 168 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_210
timestamp 1493737109
transform 1 0 212 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_233
timestamp 1493737109
transform 1 0 212 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_10
timestamp 1493737109
transform -1 0 216 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_211
timestamp 1493737109
transform 1 0 252 0 1 170
box -2 -2 2 2
use $$M3_M2  $$M3_M2_234
timestamp 1493737109
transform 1 0 252 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_212
timestamp 1493737109
transform 1 0 244 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_235
timestamp 1493737109
transform 1 0 244 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_213
timestamp 1493737109
transform 1 0 228 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_236
timestamp 1493737109
transform 1 0 228 0 1 140
box -3 -3 3 3
use FILL  FILL_25
timestamp 1493737109
transform -1 0 224 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_214
timestamp 1493737109
transform 1 0 236 0 1 137
box -2 -2 2 2
use $$M3_M2  $$M3_M2_242
timestamp 1493737109
transform 1 0 236 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_237
timestamp 1493737109
transform 1 0 292 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_215
timestamp 1493737109
transform 1 0 313 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_238
timestamp 1493737109
transform 1 0 313 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_239
timestamp 1493737109
transform 1 0 292 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_216
timestamp 1493737109
transform 1 0 276 0 1 139
box -2 -2 2 2
use $$M3_M2  $$M3_M2_240
timestamp 1493737109
transform 1 0 276 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_217
timestamp 1493737109
transform 1 0 292 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_218
timestamp 1493737109
transform 1 0 260 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_243
timestamp 1493737109
transform 1 0 268 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_244
timestamp 1493737109
transform 1 0 260 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_219
timestamp 1493737109
transform 1 0 260 0 1 118
box -2 -2 2 2
use NAND3X1  NAND3X1_10
timestamp 1493737109
transform 1 0 224 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_245
timestamp 1493737109
transform 1 0 300 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_221
timestamp 1493737109
transform 1 0 284 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_246
timestamp 1493737109
transform 1 0 268 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_247
timestamp 1493737109
transform 1 0 284 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_222
timestamp 1493737109
transform 1 0 300 0 1 111
box -2 -2 2 2
use NOR2X1  NOR2X1_11
timestamp 1493737109
transform 1 0 256 0 1 90
box -8 -3 32 105
use INVX2  INVX2_14
timestamp 1493737109
transform 1 0 280 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_241
timestamp 1493737109
transform 1 0 316 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_220
timestamp 1493737109
transform 1 0 316 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_248
timestamp 1493737109
transform 1 0 332 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_223
timestamp 1493737109
transform 1 0 340 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_249
timestamp 1493737109
transform 1 0 332 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_224
timestamp 1493737109
transform 1 0 348 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_225
timestamp 1493737109
transform 1 0 332 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_251
timestamp 1493737109
transform 1 0 324 0 1 120
box -3 -3 3 3
use NOR2X1  NOR2X1_12
timestamp 1493737109
transform 1 0 296 0 1 90
box -8 -3 32 105
use FILL  FILL_26
timestamp 1493737109
transform -1 0 328 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_226
timestamp 1493737109
transform 1 0 340 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_250
timestamp 1493737109
transform 1 0 340 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_227
timestamp 1493737109
transform 1 0 364 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_228
timestamp 1493737109
transform 1 0 380 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_252
timestamp 1493737109
transform 1 0 380 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_253
timestamp 1493737109
transform 1 0 372 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_254
timestamp 1493737109
transform 1 0 364 0 1 110
box -3 -3 3 3
use NAND3X1  NAND3X1_11
timestamp 1493737109
transform 1 0 328 0 1 90
box -8 -3 40 105
use FILL  FILL_27
timestamp 1493737109
transform -1 0 368 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_229
timestamp 1493737109
transform 1 0 388 0 1 116
box -2 -2 2 2
use $$M3_M2  $$M3_M2_262
timestamp 1493737109
transform 1 0 388 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_257
timestamp 1493737109
transform 1 0 404 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_259
timestamp 1493737109
transform 1 0 412 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_260
timestamp 1493737109
transform 1 0 404 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_255
timestamp 1493737109
transform 1 0 436 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_258
timestamp 1493737109
transform 1 0 428 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_230
timestamp 1493737109
transform 1 0 428 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_231
timestamp 1493737109
transform 1 0 404 0 1 139
box -2 -2 2 2
use $$M3_M2  $$M3_M2_261
timestamp 1493737109
transform 1 0 420 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_232
timestamp 1493737109
transform 1 0 412 0 1 125
box -2 -2 2 2
use $$M2_M1  $$M2_M1_233
timestamp 1493737109
transform 1 0 420 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_234
timestamp 1493737109
transform 1 0 396 0 1 100
box -2 -2 2 2
use INVX2  INVX2_15
timestamp 1493737109
transform 1 0 368 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_263
timestamp 1493737109
transform 1 0 412 0 1 100
box -3 -3 3 3
use NOR2X1  NOR2X1_13
timestamp 1493737109
transform 1 0 384 0 1 90
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1493737109
transform 1 0 408 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_256
timestamp 1493737109
transform 1 0 460 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_264
timestamp 1493737109
transform 1 0 444 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_235
timestamp 1493737109
transform 1 0 460 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_236
timestamp 1493737109
transform 1 0 444 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_237
timestamp 1493737109
transform 1 0 444 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_265
timestamp 1493737109
transform 1 0 444 0 1 130
box -3 -3 3 3
use FILL  FILL_28
timestamp 1493737109
transform -1 0 440 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_266
timestamp 1493737109
transform 1 0 452 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_267
timestamp 1493737109
transform 1 0 484 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_238
timestamp 1493737109
transform 1 0 484 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_239
timestamp 1493737109
transform 1 0 492 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_240
timestamp 1493737109
transform 1 0 484 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_268
timestamp 1493737109
transform 1 0 484 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_269
timestamp 1493737109
transform 1 0 492 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_241
timestamp 1493737109
transform 1 0 460 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_270
timestamp 1493737109
transform 1 0 476 0 1 100
box -3 -3 3 3
use NAND3X1  NAND3X1_12
timestamp 1493737109
transform 1 0 440 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_271
timestamp 1493737109
transform 1 0 516 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_243
timestamp 1493737109
transform 1 0 516 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_245
timestamp 1493737109
transform 1 0 508 0 1 100
box -2 -2 2 2
use NAND3X1  NAND3X1_13
timestamp 1493737109
transform 1 0 472 0 1 90
box -8 -3 40 105
use FILL  FILL_29
timestamp 1493737109
transform -1 0 512 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_242
timestamp 1493737109
transform 1 0 540 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_272
timestamp 1493737109
transform 1 0 548 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_244
timestamp 1493737109
transform 1 0 524 0 1 122
box -2 -2 2 2
use $$M2_M1  $$M2_M1_246
timestamp 1493737109
transform 1 0 548 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_247
timestamp 1493737109
transform 1 0 540 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_273
timestamp 1493737109
transform 1 0 540 0 1 110
box -3 -3 3 3
use AOI21X1  AOI21X1_2
timestamp 1493737109
transform 1 0 512 0 1 90
box -7 -3 39 105
use $$M3_M2  $$M3_M2_274
timestamp 1493737109
transform 1 0 564 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_276
timestamp 1493737109
transform 1 0 588 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_277
timestamp 1493737109
transform 1 0 572 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_248
timestamp 1493737109
transform 1 0 580 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_249
timestamp 1493737109
transform 1 0 564 0 1 111
box -2 -2 2 2
use $$M2_M1  $$M2_M1_250
timestamp 1493737109
transform 1 0 556 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_279
timestamp 1493737109
transform 1 0 564 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_278
timestamp 1493737109
transform 1 0 580 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_251
timestamp 1493737109
transform 1 0 572 0 1 100
box -2 -2 2 2
use INVX2  INVX2_16
timestamp 1493737109
transform 1 0 544 0 1 90
box -9 -3 26 105
use NOR2X1  NOR2X1_14
timestamp 1493737109
transform 1 0 560 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_275
timestamp 1493737109
transform 1 0 604 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_280
timestamp 1493737109
transform 1 0 596 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_252
timestamp 1493737109
transform 1 0 628 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_253
timestamp 1493737109
transform 1 0 612 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_281
timestamp 1493737109
transform 1 0 612 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_255
timestamp 1493737109
transform 1 0 604 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_254
timestamp 1493737109
transform 1 0 620 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_256
timestamp 1493737109
transform 1 0 596 0 1 111
box -2 -2 2 2
use FILL  FILL_30
timestamp 1493737109
transform -1 0 592 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_282
timestamp 1493737109
transform 1 0 620 0 1 90
box -3 -3 3 3
use NOR2X1  NOR2X1_15
timestamp 1493737109
transform 1 0 592 0 1 90
box -8 -3 32 105
use INVX2  INVX2_17
timestamp 1493737109
transform 1 0 616 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_283
timestamp 1493737109
transform 1 0 652 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_257
timestamp 1493737109
transform 1 0 652 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_258
timestamp 1493737109
transform 1 0 692 0 1 139
box -2 -2 2 2
use $$M3_M2  $$M3_M2_284
timestamp 1493737109
transform 1 0 692 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_261
timestamp 1493737109
transform 1 0 644 0 1 111
box -2 -2 2 2
use FILL  FILL_31
timestamp 1493737109
transform -1 0 640 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_260
timestamp 1493737109
transform 1 0 676 0 1 117
box -2 -2 2 2
use $$M2_M1  $$M2_M1_259
timestamp 1493737109
transform 1 0 684 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_285
timestamp 1493737109
transform 1 0 684 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_262
timestamp 1493737109
transform 1 0 668 0 1 100
box -2 -2 2 2
use OR2X1  OR2X1_1
timestamp 1493737109
transform 1 0 640 0 1 90
box -8 -3 40 105
use NOR2X1  NOR2X1_16
timestamp 1493737109
transform 1 0 672 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_263
timestamp 1493737109
transform 1 0 716 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_286
timestamp 1493737109
transform 1 0 716 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_288
timestamp 1493737109
transform 1 0 708 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_266
timestamp 1493737109
transform 1 0 708 0 1 121
box -2 -2 2 2
use FILL  FILL_32
timestamp 1493737109
transform -1 0 704 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_287
timestamp 1493737109
transform 1 0 732 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_264
timestamp 1493737109
transform 1 0 724 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_265
timestamp 1493737109
transform 1 0 724 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_289
timestamp 1493737109
transform 1 0 724 0 1 130
box -3 -3 3 3
use NAND2X1  NAND2X1_7
timestamp 1493737109
transform 1 0 704 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_290
timestamp 1493737109
transform 1 0 748 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_267
timestamp 1493737109
transform 1 0 748 0 1 111
box -2 -2 2 2
use $$M2_M1  $$M2_M1_268
timestamp 1493737109
transform 1 0 740 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_291
timestamp 1493737109
transform 1 0 740 0 1 90
box -3 -3 3 3
use $$M2_M1  $$M2_M1_269
timestamp 1493737109
transform 1 0 788 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_270
timestamp 1493737109
transform 1 0 772 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_271
timestamp 1493737109
transform 1 0 764 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_292
timestamp 1493737109
transform 1 0 756 0 1 90
box -3 -3 3 3
use NOR2X1  NOR2X1_17
timestamp 1493737109
transform -1 0 752 0 1 90
box -8 -3 32 105
use FILL  FILL_33
timestamp 1493737109
transform -1 0 760 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_272
timestamp 1493737109
transform 1 0 788 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_293
timestamp 1493737109
transform 1 0 788 0 1 90
box -3 -3 3 3
use OAI21X1  OAI21X1_10
timestamp 1493737109
transform 1 0 760 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_273
timestamp 1493737109
transform 1 0 828 0 1 143
box -2 -2 2 2
use $$M2_M1  $$M2_M1_274
timestamp 1493737109
transform 1 0 812 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_275
timestamp 1493737109
transform 1 0 804 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_295
timestamp 1493737109
transform 1 0 804 0 1 110
box -3 -3 3 3
use FILL  FILL_34
timestamp 1493737109
transform -1 0 800 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_294
timestamp 1493737109
transform 1 0 828 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_276
timestamp 1493737109
transform 1 0 828 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_296
timestamp 1493737109
transform 1 0 812 0 1 90
box -3 -3 3 3
use OAI21X1  OAI21X1_11
timestamp 1493737109
transform 1 0 800 0 1 90
box -8 -3 34 105
use $$M3_M2  $$M3_M2_297
timestamp 1493737109
transform 1 0 844 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_298
timestamp 1493737109
transform 1 0 852 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_277
timestamp 1493737109
transform 1 0 844 0 1 150
box -2 -2 2 2
use FILL  FILL_35
timestamp 1493737109
transform -1 0 840 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_278
timestamp 1493737109
transform 1 0 852 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_299
timestamp 1493737109
transform 1 0 852 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_280
timestamp 1493737109
transform 1 0 860 0 1 128
box -2 -2 2 2
use $$M2_M1  $$M2_M1_281
timestamp 1493737109
transform 1 0 868 0 1 119
box -2 -2 2 2
use $$M3_M2  $$M3_M2_301
timestamp 1493737109
transform 1 0 868 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_302
timestamp 1493737109
transform 1 0 860 0 1 110
box -3 -3 3 3
use NAND2X1  NAND2X1_8
timestamp 1493737109
transform -1 0 864 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_300
timestamp 1493737109
transform 1 0 884 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_279
timestamp 1493737109
transform 1 0 884 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_282
timestamp 1493737109
transform 1 0 876 0 1 100
box -2 -2 2 2
use NOR2X1  NOR2X1_18
timestamp 1493737109
transform 1 0 864 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_303
timestamp 1493737109
transform 1 0 900 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_304
timestamp 1493737109
transform 1 0 916 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_305
timestamp 1493737109
transform 1 0 908 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_306
timestamp 1493737109
transform 1 0 900 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_283
timestamp 1493737109
transform 1 0 916 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_284
timestamp 1493737109
transform 1 0 900 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_285
timestamp 1493737109
transform 1 0 908 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_307
timestamp 1493737109
transform 1 0 908 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_308
timestamp 1493737109
transform 1 0 900 0 1 90
box -3 -3 3 3
use FILL  FILL_36
timestamp 1493737109
transform -1 0 896 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_286
timestamp 1493737109
transform 1 0 924 0 1 100
box -2 -2 2 2
use NAND2X1  NAND2X1_9
timestamp 1493737109
transform 1 0 896 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_309
timestamp 1493737109
transform 1 0 932 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_287
timestamp 1493737109
transform 1 0 932 0 1 129
box -2 -2 2 2
use $$M3_M2  $$M3_M2_311
timestamp 1493737109
transform 1 0 932 0 1 100
box -3 -3 3 3
use $$M2_M1  $$M2_M1_290
timestamp 1493737109
transform 1 0 940 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_312
timestamp 1493737109
transform 1 0 940 0 1 90
box -3 -3 3 3
use INVX2  INVX2_18
timestamp 1493737109
transform -1 0 936 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_288
timestamp 1493737109
transform 1 0 956 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_310
timestamp 1493737109
transform 1 0 956 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_289
timestamp 1493737109
transform 1 0 948 0 1 121
box -2 -2 2 2
use INVX2  INVX2_19
timestamp 1493737109
transform -1 0 952 0 1 90
box -9 -3 26 105
use FILL  FILL_37
timestamp 1493737109
transform -1 0 960 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_291
timestamp 1493737109
transform 1 0 980 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_313
timestamp 1493737109
transform 1 0 980 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_292
timestamp 1493737109
transform 1 0 988 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_294
timestamp 1493737109
transform 1 0 996 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_293
timestamp 1493737109
transform 1 0 1004 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_314
timestamp 1493737109
transform 1 0 972 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_295
timestamp 1493737109
transform 1 0 972 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_316
timestamp 1493737109
transform 1 0 972 0 1 90
box -3 -3 3 3
use INVX2  INVX2_20
timestamp 1493737109
transform -1 0 976 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_315
timestamp 1493737109
transform 1 0 1004 0 1 110
box -3 -3 3 3
use NAND3X1  NAND3X1_14
timestamp 1493737109
transform -1 0 1008 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_317
timestamp 1493737109
transform 1 0 1044 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_318
timestamp 1493737109
transform 1 0 1036 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_296
timestamp 1493737109
transform 1 0 1036 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_299
timestamp 1493737109
transform 1 0 1020 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_297
timestamp 1493737109
transform 1 0 1060 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_319
timestamp 1493737109
transform 1 0 1060 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_298
timestamp 1493737109
transform 1 0 1068 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_300
timestamp 1493737109
transform 1 0 1052 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_321
timestamp 1493737109
transform 1 0 1028 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_301
timestamp 1493737109
transform 1 0 1036 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_320
timestamp 1493737109
transform 1 0 1060 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_322
timestamp 1493737109
transform 1 0 1052 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_302
timestamp 1493737109
transform 1 0 1060 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_323
timestamp 1493737109
transform 1 0 1020 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_324
timestamp 1493737109
transform 1 0 1020 0 1 100
box -3 -3 3 3
use $$M2_M1  $$M2_M1_303
timestamp 1493737109
transform 1 0 1036 0 1 100
box -2 -2 2 2
use FILL  FILL_38
timestamp 1493737109
transform -1 0 1016 0 1 90
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1493737109
transform 1 0 1016 0 1 90
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1493737109
transform 1 0 1048 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_304
timestamp 1493737109
transform 1 0 1100 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_306
timestamp 1493737109
transform 1 0 1116 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_325
timestamp 1493737109
transform 1 0 1116 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_307
timestamp 1493737109
transform 1 0 1124 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_305
timestamp 1493737109
transform 1 0 1092 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_326
timestamp 1493737109
transform 1 0 1092 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_308
timestamp 1493737109
transform 1 0 1108 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_327
timestamp 1493737109
transform 1 0 1108 0 1 110
box -3 -3 3 3
use FILL  FILL_39
timestamp 1493737109
transform -1 0 1088 0 1 90
box -8 -3 16 105
use INVX2  INVX2_21
timestamp 1493737109
transform 1 0 1088 0 1 90
box -9 -3 26 105
use NOR2X1  NOR2X1_19
timestamp 1493737109
transform 1 0 1104 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_328
timestamp 1493737109
transform 1 0 1140 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_309
timestamp 1493737109
transform 1 0 1156 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_310
timestamp 1493737109
transform 1 0 1140 0 1 140
box -2 -2 2 2
use FILL  FILL_40
timestamp 1493737109
transform -1 0 1136 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_311
timestamp 1493737109
transform 1 0 1164 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_312
timestamp 1493737109
transform 1 0 1148 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_329
timestamp 1493737109
transform 1 0 1156 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_330
timestamp 1493737109
transform 1 0 1148 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_313
timestamp 1493737109
transform 1 0 1180 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_314
timestamp 1493737109
transform 1 0 1172 0 1 100
box -2 -2 2 2
use NAND3X1  NAND3X1_17
timestamp 1493737109
transform 1 0 1136 0 1 90
box -8 -3 40 105
use INVX2  INVX2_22
timestamp 1493737109
transform -1 0 1184 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_332
timestamp 1493737109
transform 1 0 1212 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_315
timestamp 1493737109
transform 1 0 1212 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_316
timestamp 1493737109
transform 1 0 1196 0 1 140
box -2 -2 2 2
use FILL  FILL_41
timestamp 1493737109
transform -1 0 1192 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_317
timestamp 1493737109
transform 1 0 1204 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_333
timestamp 1493737109
transform 1 0 1204 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_318
timestamp 1493737109
transform 1 0 1204 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_334
timestamp 1493737109
transform 1 0 1204 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_331
timestamp 1493737109
transform 1 0 1228 0 1 170
box -3 -3 3 3
use NAND3X1  NAND3X1_18
timestamp 1493737109
transform 1 0 1192 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_335
timestamp 1493737109
transform 1 0 1252 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_319
timestamp 1493737109
transform 1 0 1252 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_320
timestamp 1493737109
transform 1 0 1236 0 1 140
box -2 -2 2 2
use FILL  FILL_42
timestamp 1493737109
transform -1 0 1232 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_321
timestamp 1493737109
transform 1 0 1244 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_336
timestamp 1493737109
transform 1 0 1244 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_337
timestamp 1493737109
transform 1 0 1244 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_338
timestamp 1493737109
transform 1 0 1284 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_340
timestamp 1493737109
transform 1 0 1276 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_322
timestamp 1493737109
transform 1 0 1276 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_339
timestamp 1493737109
transform 1 0 1300 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_324
timestamp 1493737109
transform 1 0 1284 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_323
timestamp 1493737109
transform 1 0 1292 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_341
timestamp 1493737109
transform 1 0 1284 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_325
timestamp 1493737109
transform 1 0 1284 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_342
timestamp 1493737109
transform 1 0 1292 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_343
timestamp 1493737109
transform 1 0 1284 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_326
timestamp 1493737109
transform 1 0 1252 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_344
timestamp 1493737109
transform 1 0 1268 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_345
timestamp 1493737109
transform 1 0 1252 0 1 90
box -3 -3 3 3
use $$M3_M2  $$M3_M2_346
timestamp 1493737109
transform 1 0 1268 0 1 90
box -3 -3 3 3
use NAND3X1  NAND3X1_19
timestamp 1493737109
transform 1 0 1232 0 1 90
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1493737109
transform -1 0 1296 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_347
timestamp 1493737109
transform 1 0 1324 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_348
timestamp 1493737109
transform 1 0 1316 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_349
timestamp 1493737109
transform 1 0 1324 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_327
timestamp 1493737109
transform 1 0 1324 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_350
timestamp 1493737109
transform 1 0 1308 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_328
timestamp 1493737109
transform 1 0 1308 0 1 111
box -2 -2 2 2
use FILL  FILL_43
timestamp 1493737109
transform -1 0 1304 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_329
timestamp 1493737109
transform 1 0 1324 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_351
timestamp 1493737109
transform 1 0 1324 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_331
timestamp 1493737109
transform 1 0 1332 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_353
timestamp 1493737109
transform 1 0 1324 0 1 90
box -3 -3 3 3
use INVX1  INVX1_1
timestamp 1493737109
transform 1 0 1304 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_330
timestamp 1493737109
transform 1 0 1348 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_352
timestamp 1493737109
transform 1 0 1364 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_354
timestamp 1493737109
transform 1 0 1356 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_355
timestamp 1493737109
transform 1 0 1380 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_332
timestamp 1493737109
transform 1 0 1372 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_356
timestamp 1493737109
transform 1 0 1364 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_333
timestamp 1493737109
transform 1 0 1364 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_341
timestamp 1493737109
transform 1 0 1342 0 1 90
box -2 -2 2 2
use $$M3_M2  $$M3_M2_361
timestamp 1493737109
transform 1 0 1342 0 1 90
box -3 -3 3 3
use NOR2X1  NOR2X1_20
timestamp 1493737109
transform 1 0 1320 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_362
timestamp 1493737109
transform 1 0 1356 0 1 90
box -3 -3 3 3
use FILL  FILL_44
timestamp 1493737109
transform -1 0 1352 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_334
timestamp 1493737109
transform 1 0 1388 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_357
timestamp 1493737109
transform 1 0 1412 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_335
timestamp 1493737109
transform 1 0 1420 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_358
timestamp 1493737109
transform 1 0 1420 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_336
timestamp 1493737109
transform 1 0 1428 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_337
timestamp 1493737109
transform 1 0 1412 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_339
timestamp 1493737109
transform 1 0 1404 0 1 127
box -2 -2 2 2
use $$M3_M2  $$M3_M2_359
timestamp 1493737109
transform 1 0 1396 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_340
timestamp 1493737109
transform 1 0 1372 0 1 100
box -2 -2 2 2
use INVX2  INVX2_23
timestamp 1493737109
transform -1 0 1368 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_360
timestamp 1493737109
transform 1 0 1380 0 1 100
box -3 -3 3 3
use OAI21X1  OAI21X1_12
timestamp 1493737109
transform -1 0 1400 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_338
timestamp 1493737109
transform 1 0 1420 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_363
timestamp 1493737109
transform 1 0 1420 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_369
timestamp 1493737109
transform 1 0 1412 0 1 90
box -3 -3 3 3
use FILL  FILL_45
timestamp 1493737109
transform -1 0 1408 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_370
timestamp 1493737109
transform 1 0 1428 0 1 90
box -3 -3 3 3
use NAND3X1  NAND3X1_21
timestamp 1493737109
transform 1 0 1408 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_364
timestamp 1493737109
transform 1 0 1476 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_365
timestamp 1493737109
transform 1 0 1460 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_342
timestamp 1493737109
transform 1 0 1476 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_343
timestamp 1493737109
transform 1 0 1460 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_344
timestamp 1493737109
transform 1 0 1452 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_366
timestamp 1493737109
transform 1 0 1452 0 1 110
box -3 -3 3 3
use FILL  FILL_46
timestamp 1493737109
transform -1 0 1448 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_367
timestamp 1493737109
transform 1 0 1492 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_346
timestamp 1493737109
transform 1 0 1492 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_347
timestamp 1493737109
transform 1 0 1500 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_348
timestamp 1493737109
transform 1 0 1484 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_349
timestamp 1493737109
transform 1 0 1476 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_371
timestamp 1493737109
transform 1 0 1468 0 1 90
box -3 -3 3 3
use OAI21X1  OAI21X1_13
timestamp 1493737109
transform 1 0 1448 0 1 90
box -8 -3 34 105
use $$M3_M2  $$M3_M2_372
timestamp 1493737109
transform 1 0 1484 0 1 90
box -3 -3 3 3
use INVX2  INVX2_24
timestamp 1493737109
transform 1 0 1480 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_368
timestamp 1493737109
transform 1 0 1516 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_345
timestamp 1493737109
transform 1 0 1516 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_353
timestamp 1493737109
transform 1 0 1524 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_375
timestamp 1493737109
transform 1 0 1524 0 1 130
box -3 -3 3 3
use NAND2X1  NAND2X1_10
timestamp 1493737109
transform 1 0 1496 0 1 90
box -8 -3 32 105
use FILL  FILL_47
timestamp 1493737109
transform -1 0 1528 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_373
timestamp 1493737109
transform 1 0 1540 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_374
timestamp 1493737109
transform 1 0 1548 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_350
timestamp 1493737109
transform 1 0 1540 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_351
timestamp 1493737109
transform 1 0 1556 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_352
timestamp 1493737109
transform 1 0 1548 0 1 136
box -2 -2 2 2
use $$M2_M1  $$M2_M1_354
timestamp 1493737109
transform 1 0 1540 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_376
timestamp 1493737109
transform 1 0 1540 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_377
timestamp 1493737109
transform 1 0 1556 0 1 120
box -3 -3 3 3
use NAND3X1  NAND3X1_22
timestamp 1493737109
transform -1 0 1560 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_357
timestamp 1493737109
transform 1 0 1572 0 1 121
box -2 -2 2 2
use FILL  FILL_48
timestamp 1493737109
transform -1 0 1568 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_355
timestamp 1493737109
transform 1 0 1580 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_378
timestamp 1493737109
transform 1 0 1588 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_379
timestamp 1493737109
transform 1 0 1588 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_356
timestamp 1493737109
transform 1 0 1588 0 1 127
box -2 -2 2 2
use INVX2  INVX2_25
timestamp 1493737109
transform 1 0 1568 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_358
timestamp 1493737109
transform 1 0 1596 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_359
timestamp 1493737109
transform 1 0 1604 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_360
timestamp 1493737109
transform 1 0 1604 0 1 130
box -2 -2 2 2
use INVX2  INVX2_26
timestamp 1493737109
transform 1 0 1584 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_380
timestamp 1493737109
transform 1 0 1628 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_361
timestamp 1493737109
transform 1 0 1620 0 1 117
box -2 -2 2 2
use NOR2X1  NOR2X1_21
timestamp 1493737109
transform -1 0 1624 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_362
timestamp 1493737109
transform 1 0 1652 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_381
timestamp 1493737109
transform 1 0 1644 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_363
timestamp 1493737109
transform 1 0 1644 0 1 127
box -2 -2 2 2
use $$M3_M2  $$M3_M2_384
timestamp 1493737109
transform 1 0 1652 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_367
timestamp 1493737109
transform 1 0 1636 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_385
timestamp 1493737109
transform 1 0 1636 0 1 100
box -3 -3 3 3
use FILL  FILL_49
timestamp 1493737109
transform -1 0 1632 0 1 90
box -8 -3 16 105
use INVX2  INVX2_27
timestamp 1493737109
transform -1 0 1648 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_383
timestamp 1493737109
transform 1 0 1668 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_366
timestamp 1493737109
transform 1 0 1660 0 1 123
box -2 -2 2 2
use INVX2  INVX2_28
timestamp 1493737109
transform -1 0 1664 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_364
timestamp 1493737109
transform 1 0 1684 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_382
timestamp 1493737109
transform 1 0 1692 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_365
timestamp 1493737109
transform 1 0 1692 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_368
timestamp 1493737109
transform 1 0 1676 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_386
timestamp 1493737109
transform 1 0 1684 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_369
timestamp 1493737109
transform 1 0 1692 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_387
timestamp 1493737109
transform 1 0 1716 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_389
timestamp 1493737109
transform 1 0 1676 0 1 120
box -3 -3 3 3
use FILL  FILL_50
timestamp 1493737109
transform -1 0 1672 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_372
timestamp 1493737109
transform 1 0 1708 0 1 127
box -2 -2 2 2
use NAND3X1  NAND3X1_23
timestamp 1493737109
transform 1 0 1672 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_370
timestamp 1493737109
transform 1 0 1724 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_371
timestamp 1493737109
transform 1 0 1732 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_388
timestamp 1493737109
transform 1 0 1732 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_373
timestamp 1493737109
transform 1 0 1732 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_390
timestamp 1493737109
transform 1 0 1724 0 1 100
box -3 -3 3 3
use NAND2X1  NAND2X1_11
timestamp 1493737109
transform 1 0 1704 0 1 90
box -8 -3 32 105
use FILL  FILL_51
timestamp 1493737109
transform -1 0 1736 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_374
timestamp 1493737109
transform 1 0 1750 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_391
timestamp 1493737109
transform 1 0 1764 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_375
timestamp 1493737109
transform 1 0 1756 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_376
timestamp 1493737109
transform 1 0 1764 0 1 124
box -2 -2 2 2
use OAI21X1  OAI21X1_14
timestamp 1493737109
transform -1 0 1768 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_377
timestamp 1493737109
transform 1 0 1788 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_392
timestamp 1493737109
transform 1 0 1788 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_378
timestamp 1493737109
transform 1 0 1828 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_380
timestamp 1493737109
transform 1 0 1804 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_381
timestamp 1493737109
transform 1 0 1796 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_393
timestamp 1493737109
transform 1 0 1828 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_379
timestamp 1493737109
transform 1 0 1852 0 1 143
box -2 -2 2 2
use $$M2_M1  $$M2_M1_382
timestamp 1493737109
transform 1 0 1836 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_394
timestamp 1493737109
transform 1 0 1836 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_395
timestamp 1493737109
transform 1 0 1804 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_384
timestamp 1493737109
transform 1 0 1828 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_385
timestamp 1493737109
transform 1 0 1786 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_396
timestamp 1493737109
transform 1 0 1786 0 1 100
box -3 -3 3 3
use $$M2_M1  $$M2_M1_386
timestamp 1493737109
transform 1 0 1812 0 1 100
box -2 -2 2 2
use FILL  FILL_52
timestamp 1493737109
transform -1 0 1776 0 1 90
box -8 -3 16 105
use NAND3X1  NAND3X1_24
timestamp 1493737109
transform -1 0 1808 0 1 90
box -8 -3 40 105
use INVX2  INVX2_29
timestamp 1493737109
transform -1 0 1824 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_383
timestamp 1493737109
transform 1 0 1844 0 1 124
box -2 -2 2 2
use $$M3_M2  $$M3_M2_397
timestamp 1493737109
transform 1 0 1844 0 1 120
box -3 -3 3 3
use NAND2X1  NAND2X1_12
timestamp 1493737109
transform -1 0 1848 0 1 90
box -8 -3 32 105
use FILL  FILL_53
timestamp 1493737109
transform -1 0 1856 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_387
timestamp 1493737109
transform 1 0 1870 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_390
timestamp 1493737109
transform 1 0 1876 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_399
timestamp 1493737109
transform 1 0 1876 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_388
timestamp 1493737109
transform 1 0 1903 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_398
timestamp 1493737109
transform 1 0 1903 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_389
timestamp 1493737109
transform 1 0 1892 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_391
timestamp 1493737109
transform 1 0 1884 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_400
timestamp 1493737109
transform 1 0 1884 0 1 110
box -3 -3 3 3
use OAI21X1  OAI21X1_15
timestamp 1493737109
transform -1 0 1888 0 1 90
box -8 -3 34 105
use FILL  FILL_54
timestamp 1493737109
transform -1 0 1896 0 1 90
box -8 -3 16 105
use NOR2X1  NOR2X1_22
timestamp 1493737109
transform -1 0 1920 0 1 90
box -8 -3 32 105
use FILL  FILL_55
timestamp 1493737109
transform -1 0 1928 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_392
timestamp 1493737109
transform 1 0 1996 0 1 136
box -2 -2 2 2
use $$M2_M1  $$M2_M1_393
timestamp 1493737109
transform 1 0 2004 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_394
timestamp 1493737109
transform 1 0 1940 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_401
timestamp 1493737109
transform 1 0 1940 0 1 110
box -3 -3 3 3
use FILL  FILL_56
timestamp 1493737109
transform -1 0 1936 0 1 90
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_3
timestamp 1493737109
transform -1 0 2032 0 1 90
box -8 -3 104 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1493737109
transform 1 0 2049 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1493737109
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_402
timestamp 1493737109
transform 1 0 460 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_403
timestamp 1493737109
transform 1 0 524 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_404
timestamp 1493737109
transform 1 0 644 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_405
timestamp 1493737109
transform 1 0 748 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_406
timestamp 1493737109
transform 1 0 764 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_407
timestamp 1493737109
transform 1 0 844 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_408
timestamp 1493737109
transform 1 0 924 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_409
timestamp 1493737109
transform 1 0 948 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_410
timestamp 1493737109
transform 1 0 1028 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_411
timestamp 1493737109
transform 1 0 1180 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_412
timestamp 1493737109
transform 1 0 1324 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_413
timestamp 1493737109
transform 1 0 1364 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_414
timestamp 1493737109
transform 1 0 1460 0 1 80
box -3 -3 3 3
use $$M3_M2  $$M3_M2_415
timestamp 1493737109
transform 1 0 700 0 1 70
box -3 -3 3 3
use $$M3_M2  $$M3_M2_416
timestamp 1493737109
transform 1 0 1020 0 1 70
box -3 -3 3 3
use $$M3_M2  $$M3_M2_417
timestamp 1493737109
transform 1 0 1132 0 1 70
box -3 -3 3 3
use $$M3_M2  $$M3_M2_418
timestamp 1493737109
transform 1 0 1316 0 1 70
box -3 -3 3 3
use $$M3_M2_1500_1500_1_2  $$M3_M2_1500_1500_1_2_2
timestamp 1493737109
transform 1 0 1342 0 1 72
box -3 -6 3 5
use $$M3_M2  $$M3_M2_419
timestamp 1493737109
transform 1 0 1364 0 1 70
box -3 -3 3 3
use $$M3_M2  $$M3_M2_420
timestamp 1493737109
transform 1 0 1812 0 1 70
box -3 -3 3 3
use $$M2_M1_1500_1500_1_3  $$M2_M1_1500_1500_1_3_2
timestamp 1493737109
transform 1 0 1342 0 1 72
box -2 -7 2 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1493737109
transform 1 0 2049 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_421
timestamp 1493737109
transform 1 0 500 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_422
timestamp 1493737109
transform 1 0 1124 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_423
timestamp 1493737109
transform 1 0 1252 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_424
timestamp 1493737109
transform 1 0 1356 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_425
timestamp 1493737109
transform 1 0 1436 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1493737109
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M3_M2  $$M3_M2_426
timestamp 1493737109
transform 1 0 332 0 1 50
box -3 -3 3 3
use $$M3_M2  $$M3_M2_427
timestamp 1493737109
transform 1 0 876 0 1 50
box -3 -3 3 3
use $$M3_M2  $$M3_M2_428
timestamp 1493737109
transform 1 0 1028 0 1 50
box -3 -3 3 3
use $$M3_M2  $$M3_M2_429
timestamp 1493737109
transform 1 0 1324 0 1 50
box -3 -3 3 3
use $$M3_M2  $$M3_M2_432
timestamp 1493737109
transform 1 0 772 0 1 40
box -3 -3 3 3
use $$M3_M2  $$M3_M2_433
timestamp 1493737109
transform 1 0 828 0 1 40
box -3 -3 3 3
use $$M3_M2  $$M3_M2_434
timestamp 1493737109
transform 1 0 1084 0 1 40
box -3 -3 3 3
use $$M3_M2  $$M3_M2_435
timestamp 1493737109
transform 1 0 1100 0 1 40
box -3 -3 3 3
use $$M3_M2_1500_1500_1_2  $$M3_M2_1500_1500_1_2_3
timestamp 1493737109
transform 1 0 1333 0 1 47
box -3 -6 3 5
use $$M3_M2  $$M3_M2_430
timestamp 1493737109
transform 1 0 1348 0 1 50
box -3 -3 3 3
use $$M3_M2  $$M3_M2_431
timestamp 1493737109
transform 1 0 1724 0 1 50
box -3 -3 3 3
use $$M2_M1_1500_1500_1_3  $$M2_M1_1500_1500_1_3_3
timestamp 1493737109
transform 1 0 1333 0 1 47
box -2 -7 2 7
use $$M3_M2  $$M3_M2_436
timestamp 1493737109
transform 1 0 1476 0 1 40
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1493737109
transform 1 0 2074 0 1 47
box -7 -7 7 7
use $$M2_M1  $$M2_M1_395
timestamp 1493737109
transform 1 0 44 0 1 30
box -2 -2 2 2
use $$M3_M2  $$M3_M2_437
timestamp 1493737109
transform 1 0 300 0 1 30
box -3 -3 3 3
use $$M3_M2  $$M3_M2_438
timestamp 1493737109
transform 1 0 396 0 1 30
box -3 -3 3 3
use $$M3_M2  $$M3_M2_439
timestamp 1493737109
transform 1 0 436 0 1 30
box -3 -3 3 3
use $$M2_M1  $$M2_M1_396
timestamp 1493737109
transform 1 0 756 0 1 30
box -2 -2 2 2
use $$M2_M1  $$M2_M1_397
timestamp 1493737109
transform 1 0 860 0 1 30
box -2 -2 2 2
use $$M3_M2  $$M3_M2_440
timestamp 1493737109
transform 1 0 1004 0 1 30
box -3 -3 3 3
use $$M3_M2  $$M3_M2_441
timestamp 1493737109
transform 1 0 1284 0 1 30
box -3 -3 3 3
use $$M3_M2  $$M3_M2_442
timestamp 1493737109
transform 1 0 1436 0 1 30
box -3 -3 3 3
use $$M2_M1  $$M2_M1_398
timestamp 1493737109
transform 1 0 1452 0 1 30
box -2 -2 2 2
use $$M2_M1  $$M2_M1_399
timestamp 1493737109
transform 1 0 1460 0 1 30
box -2 -2 2 2
use $$M2_M1  $$M2_M1_400
timestamp 1493737109
transform 1 0 1796 0 1 30
box -2 -2 2 2
use $$M3_M2  $$M3_M2_443
timestamp 1493737109
transform 1 0 1836 0 1 30
box -3 -3 3 3
use $$M3_M2  $$M3_M2_444
timestamp 1493737109
transform 1 0 508 0 1 20
box -3 -3 3 3
use $$M2_M1  $$M2_M1_401
timestamp 1493737109
transform 1 0 604 0 1 20
box -2 -2 2 2
use $$M2_M1  $$M2_M1_402
timestamp 1493737109
transform 1 0 1140 0 1 20
box -2 -2 2 2
use $$M2_M1  $$M2_M1_403
timestamp 1493737109
transform 1 0 1220 0 1 20
box -2 -2 2 2
use $$M2_M1  $$M2_M1_404
timestamp 1493737109
transform 1 0 1572 0 1 20
box -2 -2 2 2
use $$M3_M2  $$M3_M2_445
timestamp 1493737109
transform 1 0 1852 0 1 20
box -3 -3 3 3
use $$M2_M1  $$M2_M1_405
timestamp 1493737109
transform 1 0 404 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_446
timestamp 1493737109
transform 1 0 548 0 1 10
box -3 -3 3 3
use $$M2_M1  $$M2_M1_406
timestamp 1493737109
transform 1 0 596 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_447
timestamp 1493737109
transform 1 0 804 0 1 10
box -3 -3 3 3
use $$M2_M1  $$M2_M1_407
timestamp 1493737109
transform 1 0 916 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_448
timestamp 1493737109
transform 1 0 932 0 1 10
box -3 -3 3 3
use $$M3_M2  $$M3_M2_449
timestamp 1493737109
transform 1 0 1012 0 1 10
box -3 -3 3 3
use $$M3_M2  $$M3_M2_450
timestamp 1493737109
transform 1 0 1036 0 1 10
box -3 -3 3 3
use $$M2_M1  $$M2_M1_408
timestamp 1493737109
transform 1 0 1172 0 1 10
box -2 -2 2 2
use $$M2_M1  $$M2_M1_409
timestamp 1493737109
transform 1 0 1252 0 1 10
box -2 -2 2 2
use $$M2_M1  $$M2_M1_410
timestamp 1493737109
transform 1 0 1308 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_451
timestamp 1493737109
transform 1 0 1372 0 1 10
box -3 -3 3 3
use $$M3_M2  $$M3_M2_452
timestamp 1493737109
transform 1 0 1412 0 1 10
box -3 -3 3 3
use $$M2_M1  $$M2_M1_411
timestamp 1493737109
transform 1 0 1444 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_453
timestamp 1493737109
transform 1 0 1460 0 1 10
box -3 -3 3 3
use $$M2_M1  $$M2_M1_412
timestamp 1493737109
transform 1 0 1468 0 1 10
box -2 -2 2 2
use $$M3_M2  $$M3_M2_454
timestamp 1493737109
transform 1 0 68 0 1 3
box -3 -3 3 3
<< labels >>
flabel metal3 2 320 2 320 4 FreeSans 26 0 0 0 clk
flabel metal2 44 378 44 378 4 FreeSans 26 0 0 0 reset
flabel metal2 1332 378 1332 378 4 FreeSans 26 0 0 0 memwrite
flabel metal2 636 1 636 1 4 FreeSans 26 0 0 0 regdst
flabel metal2 404 1 404 1 4 FreeSans 26 0 0 0 memtoreg
flabel metal2 132 1 132 1 4 FreeSans 26 0 0 0 op[4]
flabel metal2 268 1 268 1 4 FreeSans 26 0 0 0 op[0]
flabel metal2 500 1 500 1 4 FreeSans 26 0 0 0 funct[3]
flabel metal2 868 1 868 1 4 FreeSans 26 0 0 0 pcsrc[0]
flabel metal2 436 1 436 1 4 FreeSans 26 0 0 0 funct[5]
flabel metal2 572 1 572 1 4 FreeSans 26 0 0 0 funct[1]
flabel metal2 236 1 236 1 4 FreeSans 26 0 0 0 op[1]
flabel metal2 204 1 204 1 4 FreeSans 26 0 0 0 op[2]
flabel metal2 68 1 68 1 4 FreeSans 26 0 0 0 irwrite[3]
flabel metal2 532 1 532 1 4 FreeSans 26 0 0 0 funct[2]
flabel metal2 172 1 172 1 4 FreeSans 26 0 0 0 op[3]
flabel metal2 604 1 604 1 4 FreeSans 26 0 0 0 funct[0]
flabel metal2 804 1 804 1 4 FreeSans 26 0 0 0 alusrcb[1]
flabel metal2 900 1 900 1 4 FreeSans 26 0 0 0 pcsrc[1]
flabel metal2 468 1 468 1 4 FreeSans 26 0 0 0 funct[4]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 iord
flabel metal2 300 1 300 1 4 FreeSans 26 0 0 0 irwrite[2]
flabel metal2 100 1 100 1 4 FreeSans 26 0 0 0 op[5]
flabel metal2 332 1 332 1 4 FreeSans 26 0 0 0 irwrite[1]
flabel metal2 1132 1 1132 1 4 FreeSans 26 0 0 0 zero
flabel metal2 372 1 372 1 4 FreeSans 26 0 0 0 irwrite[0]
flabel metal2 932 1 932 1 4 FreeSans 26 0 0 0 pcen
flabel metal2 668 1 668 1 4 FreeSans 26 0 0 0 regwrite
flabel metal2 1068 1 1068 1 4 FreeSans 26 0 0 0 alucontrol[0]
flabel metal2 1100 1 1100 1 4 FreeSans 26 0 0 0 alucontrol[1]
flabel metal2 700 1 700 1 4 FreeSans 26 0 0 0 alucontrol[2]
flabel metal2 732 1 732 1 4 FreeSans 26 0 0 0 alucontrol[3]
flabel metal2 1036 1 1036 1 4 FreeSans 26 0 0 0 alucontrol[4]
flabel metal2 1004 1 1004 1 4 FreeSans 26 0 0 0 alucontrol[5]
flabel metal2 972 1 972 1 4 FreeSans 26 0 0 0 alucontrol[6]
flabel metal2 836 1 836 1 4 FreeSans 26 0 0 0 alusrca
flabel metal2 772 1 772 1 4 FreeSans 26 0 0 0 alusrcb[0]
<< end >>
