magic
tech scmos
timestamp 1490995571
<< m2contact >>
rect -2 -2 2 2
<< end >>
