magic
tech scmos
timestamp 1494182186
<< metal1 >>
rect 3919 3799 4004 3895
rect 3716 3441 3919 3444
rect 3716 3432 3855 3441
rect 3716 3429 3919 3432
rect 3698 3416 3991 3419
rect 3698 3407 3927 3416
rect 3698 3404 3991 3407
rect 1285 2515 1287 2517
rect 3300 2513 3302 2515
rect 1285 2405 1287 2407
rect 3300 2403 3302 2405
rect 1285 2295 1287 2297
rect 3300 2293 3302 2295
rect 1285 2185 1287 2187
rect 3300 2183 3302 2185
rect 1285 2074 1287 2076
rect 3300 2073 3302 2075
rect 1285 1965 1287 1967
rect 3300 1963 3302 1965
rect 1285 1855 1287 1857
rect 3300 1853 3302 1855
rect 1285 1745 1287 1747
rect 3298 1743 3300 1745
<< m2contact >>
rect 3855 3799 3919 3895
rect 3855 3432 3919 3441
rect 3927 3407 3991 3416
<< metal2 >>
rect 1034 3993 1038 3994
rect 998 3959 1008 3963
rect 1004 3921 1008 3959
rect 1004 3916 1008 3917
rect 1006 2222 1010 2459
rect 1013 2332 1017 2759
rect 1020 2442 1024 3059
rect 1027 2552 1031 3359
rect 1027 2547 1031 2548
rect 1020 2437 1024 2438
rect 1013 2327 1017 2328
rect 1006 2163 1010 2164
rect 1006 2112 1010 2159
rect 1020 2002 1024 2003
rect 1013 1892 1017 1893
rect 1006 1782 1010 1783
rect 1006 1050 1010 1778
rect 1013 1350 1017 1888
rect 1020 1863 1024 1998
rect 1034 1762 1038 3989
rect 1041 3984 1045 3985
rect 1041 1872 1045 3980
rect 1048 3975 1052 3976
rect 1048 1982 1052 3971
rect 1055 3966 1059 3967
rect 1055 2092 1059 3962
rect 1062 3957 1066 3958
rect 1062 2202 1066 3953
rect 1069 3948 1073 3949
rect 1069 2312 1073 3944
rect 1076 3939 1080 3940
rect 1076 2422 1080 3935
rect 1083 3930 1087 3931
rect 1083 2532 1087 3926
rect 1259 3922 1263 4004
rect 1346 3993 1350 4002
rect 1346 3988 1350 3989
rect 1646 3984 1650 4002
rect 1646 3979 1650 3980
rect 1946 3975 1950 4002
rect 1946 3970 1950 3971
rect 2246 3966 2250 4002
rect 2246 3961 2250 3962
rect 2546 3957 2550 4002
rect 2546 3952 2550 3953
rect 2846 3948 2850 4002
rect 2846 3943 2850 3944
rect 2984 3993 2988 3994
rect 1259 3918 1267 3922
rect 1263 3484 1267 3918
rect 1279 3921 1283 3922
rect 1263 3007 1267 3480
rect 1271 3663 1275 3664
rect 1271 3426 1275 3659
rect 1271 3007 1275 3422
rect 1279 3008 1283 3917
rect 2984 3483 2988 3989
rect 3146 3939 3150 4002
rect 3146 3934 3150 3935
rect 3446 3930 3450 4002
rect 3746 3993 3750 4002
rect 3746 3988 3750 3989
rect 3446 3925 3450 3926
rect 3855 3441 3919 3799
rect 1697 3113 1699 3115
rect 3855 3027 3919 3432
rect 3927 3500 4006 3596
rect 3927 3416 3991 3500
rect 3927 3043 3991 3407
rect 3216 3005 3218 3007
rect 3248 3005 3250 3007
rect 3304 2570 3306 2572
rect 1083 2527 1087 2528
rect 2191 2542 2195 2543
rect 1076 2417 1080 2418
rect 2183 2432 2187 2433
rect 1069 2307 1073 2308
rect 2175 2322 2179 2323
rect 1062 2197 1066 2198
rect 1623 2212 1627 2213
rect 1055 2087 1059 2088
rect 1463 2102 1467 2103
rect 1048 1977 1052 1978
rect 1455 1992 1459 1993
rect 1041 1867 1045 1868
rect 1447 1882 1451 1883
rect 1034 1757 1038 1758
rect 1439 1772 1443 1773
rect 1250 1020 1254 1021
rect 1250 998 1254 1016
rect 1439 1020 1443 1768
rect 1439 1015 1443 1016
rect 1447 1011 1451 1878
rect 1455 1020 1459 1988
rect 1463 1029 1467 2098
rect 1623 1038 1627 2208
rect 2175 1047 2179 2318
rect 2183 1056 2187 2428
rect 2191 1065 2195 2538
rect 2191 1060 2195 1061
rect 3350 1065 3354 1066
rect 2183 1051 2187 1052
rect 3050 1056 3054 1057
rect 2175 1042 2179 1043
rect 2750 1047 2754 1048
rect 1623 1033 1627 1034
rect 1463 1024 1467 1025
rect 2150 1029 2154 1030
rect 1455 1015 1459 1016
rect 1850 1020 1854 1021
rect 1447 999 1451 1007
rect 1550 1011 1554 1012
rect 1550 991 1554 1007
rect 1850 998 1854 1016
rect 2150 1000 2154 1025
rect 2150 998 2155 1000
rect 2450 998 2454 1034
rect 2750 998 2754 1043
rect 3050 998 3054 1052
rect 3350 1000 3354 1061
rect 3350 998 3355 1000
<< m3contact >>
rect 1034 3989 1038 3993
rect 1004 3917 1008 3921
rect 998 3659 1002 3663
rect 998 3359 1002 3363
rect 1027 3359 1031 3363
rect 998 3059 1002 3063
rect 1020 3059 1024 3063
rect 998 2759 1002 2763
rect 1013 2759 1017 2763
rect 998 2459 1002 2463
rect 1006 2459 1010 2463
rect 1027 2548 1031 2552
rect 1020 2438 1024 2442
rect 1013 2328 1017 2332
rect 1006 2218 1010 2222
rect 998 2159 1002 2163
rect 1006 2159 1010 2163
rect 1006 2108 1010 2112
rect 1020 1998 1024 2002
rect 1013 1888 1017 1892
rect 998 1859 1002 1863
rect 1006 1778 1010 1782
rect 998 1346 1002 1350
rect 1020 1859 1024 1863
rect 1041 3980 1045 3984
rect 1048 3971 1052 3975
rect 1055 3962 1059 3966
rect 1062 3953 1066 3957
rect 1069 3944 1073 3948
rect 1076 3935 1080 3939
rect 1083 3926 1087 3930
rect 1346 3989 1350 3993
rect 1646 3980 1650 3984
rect 1946 3971 1950 3975
rect 2246 3962 2250 3966
rect 2546 3953 2550 3957
rect 2846 3944 2850 3948
rect 2984 3989 2988 3993
rect 1279 3917 1283 3921
rect 1263 3480 1267 3484
rect 1271 3659 1275 3663
rect 1271 3422 1275 3426
rect 1673 3480 1677 3484
rect 3146 3935 3150 3939
rect 3746 3989 3750 3993
rect 3446 3926 3450 3930
rect 1083 2528 1087 2532
rect 2191 2538 2195 2542
rect 1076 2418 1080 2422
rect 2183 2428 2187 2432
rect 1069 2308 1073 2312
rect 2175 2318 2179 2322
rect 1062 2198 1066 2202
rect 1623 2208 1627 2212
rect 1055 2088 1059 2092
rect 1463 2098 1467 2102
rect 1048 1978 1052 1982
rect 1455 1988 1459 1992
rect 1041 1868 1045 1872
rect 1447 1878 1451 1882
rect 1034 1758 1038 1762
rect 1439 1768 1443 1772
rect 1013 1346 1017 1350
rect 998 1046 1002 1050
rect 1006 1046 1010 1050
rect 1250 1016 1254 1020
rect 1439 1016 1443 1020
rect 2191 1061 2195 1065
rect 3350 1061 3354 1065
rect 2183 1052 2187 1056
rect 3050 1052 3054 1056
rect 2175 1043 2179 1047
rect 2750 1043 2754 1047
rect 1623 1034 1627 1038
rect 2450 1034 2454 1038
rect 1463 1025 1467 1029
rect 2150 1025 2154 1029
rect 1455 1016 1459 1020
rect 1850 1016 1854 1020
rect 1447 1007 1451 1011
rect 1550 1007 1554 1011
<< metal3 >>
rect 1033 3993 1351 3994
rect 1033 3989 1034 3993
rect 1038 3989 1346 3993
rect 1350 3989 1351 3993
rect 1033 3988 1351 3989
rect 2983 3993 3751 3994
rect 2983 3989 2984 3993
rect 2988 3989 3746 3993
rect 3750 3989 3751 3993
rect 2983 3988 3751 3989
rect 1040 3984 1651 3985
rect 1040 3980 1041 3984
rect 1045 3980 1646 3984
rect 1650 3980 1651 3984
rect 1040 3979 1651 3980
rect 1047 3975 1951 3976
rect 1047 3971 1048 3975
rect 1052 3971 1946 3975
rect 1950 3971 1951 3975
rect 1047 3970 1951 3971
rect 1054 3966 2251 3967
rect 1054 3962 1055 3966
rect 1059 3962 2246 3966
rect 2250 3962 2251 3966
rect 1054 3961 2251 3962
rect 1061 3957 2551 3958
rect 1061 3953 1062 3957
rect 1066 3953 2546 3957
rect 2550 3953 2551 3957
rect 1061 3952 2551 3953
rect 1068 3948 2851 3949
rect 1068 3944 1069 3948
rect 1073 3944 2846 3948
rect 2850 3944 2851 3948
rect 1068 3943 2851 3944
rect 1075 3939 3151 3940
rect 1075 3935 1076 3939
rect 1080 3935 3146 3939
rect 3150 3935 3151 3939
rect 1075 3934 3151 3935
rect 1082 3930 3451 3931
rect 1082 3926 1083 3930
rect 1087 3926 3446 3930
rect 3450 3926 3451 3930
rect 1082 3925 3451 3926
rect 1003 3921 1284 3922
rect 1003 3917 1004 3921
rect 1008 3917 1279 3921
rect 1283 3917 1284 3921
rect 1003 3916 1284 3917
rect 997 3663 1276 3664
rect 997 3659 998 3663
rect 1002 3659 1271 3663
rect 1275 3659 1276 3663
rect 997 3658 1276 3659
rect 1262 3484 1678 3485
rect 1262 3480 1263 3484
rect 1267 3480 1673 3484
rect 1677 3480 1678 3484
rect 1262 3479 1678 3480
rect 1270 3426 1662 3427
rect 1270 3422 1271 3426
rect 1275 3422 1662 3426
rect 1270 3421 1662 3422
rect 997 3363 1032 3364
rect 997 3359 998 3363
rect 1002 3359 1027 3363
rect 1031 3359 1032 3363
rect 997 3358 1032 3359
rect 997 3063 1025 3064
rect 997 3059 998 3063
rect 1002 3059 1020 3063
rect 1024 3059 1025 3063
rect 997 3058 1025 3059
rect 997 2763 1018 2764
rect 997 2759 998 2763
rect 1002 2759 1013 2763
rect 1017 2759 1018 2763
rect 997 2758 1018 2759
rect 1026 2552 1244 2553
rect 1026 2548 1027 2552
rect 1031 2548 1244 2552
rect 1026 2547 1244 2548
rect 1082 2532 1238 2533
rect 1082 2528 1083 2532
rect 1087 2528 1238 2532
rect 1971 2529 1973 2531
rect 1082 2527 1238 2528
rect 1260 2507 1262 2509
rect 3825 2507 3827 2509
rect 997 2463 1011 2464
rect 997 2459 998 2463
rect 1002 2459 1006 2463
rect 1010 2459 1011 2463
rect 997 2458 1011 2459
rect 1019 2442 1243 2443
rect 1019 2438 1020 2442
rect 1024 2438 1243 2442
rect 1019 2437 1243 2438
rect 1075 2422 1240 2423
rect 1075 2418 1076 2422
rect 1080 2418 1240 2422
rect 1972 2419 1974 2421
rect 1075 2417 1240 2418
rect 1260 2397 1262 2399
rect 3816 2396 3818 2398
rect 1012 2332 1244 2333
rect 1012 2328 1013 2332
rect 1017 2328 1244 2332
rect 1012 2327 1244 2328
rect 1068 2312 1239 2313
rect 1068 2308 1069 2312
rect 1073 2308 1239 2312
rect 1972 2308 1974 2310
rect 1068 2307 1239 2308
rect 1260 2288 1262 2290
rect 3813 2276 3815 2278
rect 1005 2222 1244 2223
rect 1005 2218 1006 2222
rect 1010 2218 1244 2222
rect 1005 2217 1244 2218
rect 1061 2202 1239 2203
rect 1061 2198 1062 2202
rect 1066 2198 1239 2202
rect 1972 2198 1974 2200
rect 1061 2197 1239 2198
rect 1260 2177 1262 2179
rect 3813 2166 3816 2168
rect 997 2163 1011 2164
rect 997 2159 998 2163
rect 1002 2159 1006 2163
rect 1010 2159 1011 2163
rect 997 2158 1011 2159
rect 1005 2112 1244 2113
rect 1005 2108 1006 2112
rect 1010 2108 1244 2112
rect 1005 2107 1244 2108
rect 1054 2092 1240 2093
rect 1054 2088 1055 2092
rect 1059 2088 1240 2092
rect 1972 2088 1974 2090
rect 1054 2087 1240 2088
rect 1260 2067 1262 2069
rect 3816 2049 3818 2051
rect 1019 2002 1243 2003
rect 1019 1998 1020 2002
rect 1024 1998 1243 2002
rect 1019 1997 1243 1998
rect 1047 1982 1240 1983
rect 1047 1978 1048 1982
rect 1052 1978 1240 1982
rect 1972 1979 1974 1981
rect 1047 1977 1240 1978
rect 1260 1958 1262 1960
rect 3814 1956 3816 1958
rect 1012 1892 1243 1893
rect 1012 1888 1013 1892
rect 1017 1888 1243 1892
rect 1012 1887 1243 1888
rect 1040 1872 1238 1873
rect 1040 1868 1041 1872
rect 1045 1868 1238 1872
rect 1972 1868 1974 1870
rect 1040 1867 1238 1868
rect 997 1863 1025 1864
rect 997 1859 998 1863
rect 1002 1859 1020 1863
rect 1024 1859 1025 1863
rect 997 1858 1025 1859
rect 1260 1848 1263 1850
rect 3815 1834 3819 1837
rect 1005 1782 1243 1783
rect 1005 1778 1006 1782
rect 1010 1778 1243 1782
rect 1005 1777 1243 1778
rect 1033 1762 1239 1763
rect 1033 1758 1034 1762
rect 1038 1758 1239 1762
rect 1973 1759 1975 1761
rect 1033 1757 1239 1758
rect 1260 1737 1262 1740
rect 3812 1737 3814 1739
rect 997 1350 1018 1351
rect 997 1346 998 1350
rect 1002 1346 1013 1350
rect 1017 1346 1018 1350
rect 997 1345 1018 1346
rect 2190 1065 3355 1066
rect 2190 1061 2191 1065
rect 2195 1061 3350 1065
rect 3354 1061 3355 1065
rect 2190 1060 3355 1061
rect 2182 1056 3055 1057
rect 2182 1052 2183 1056
rect 2187 1052 3050 1056
rect 3054 1052 3055 1056
rect 2182 1051 3055 1052
rect 997 1050 1011 1051
rect 997 1046 998 1050
rect 1002 1046 1006 1050
rect 1010 1046 1011 1050
rect 997 1045 1011 1046
rect 2174 1047 2755 1048
rect 2174 1043 2175 1047
rect 2179 1043 2750 1047
rect 2754 1043 2755 1047
rect 2174 1042 2755 1043
rect 1622 1038 2455 1039
rect 1622 1034 1623 1038
rect 1627 1034 2450 1038
rect 2454 1034 2455 1038
rect 1622 1033 2455 1034
rect 1462 1029 2155 1030
rect 1462 1025 1463 1029
rect 1467 1025 2150 1029
rect 2154 1025 2155 1029
rect 1462 1024 2155 1025
rect 1249 1020 1444 1021
rect 1249 1016 1250 1020
rect 1254 1016 1439 1020
rect 1443 1016 1444 1020
rect 1249 1015 1444 1016
rect 1454 1020 1855 1021
rect 1454 1016 1455 1020
rect 1459 1016 1850 1020
rect 1854 1016 1855 1020
rect 1454 1015 1855 1016
rect 1446 1011 1481 1012
rect 1446 1007 1447 1011
rect 1451 1007 1481 1011
rect 1446 1006 1481 1007
rect 1521 1011 1555 1012
rect 1521 1007 1550 1011
rect 1554 1007 1555 1011
rect 1521 1006 1555 1007
use alt_mips  alt_mips_0
timestamp 1494181132
transform 1 0 1115 0 1 1152
box 0 0 2876 2332
use PadFrame17  PadFrame17_0
timestamp 1491676833
transform 1 0 0 0 1 0
box 0 0 5000 5000
<< labels >>
rlabel space 3702 3437 3702 3437 1 Vdd!
rlabel space 3682 3412 3682 3412 1 Gnd!
rlabel metal2 3351 1007 3351 1007 1 writedata7
rlabel metal2 3051 1008 3051 1008 1 writedata6
rlabel metal2 2752 1007 2752 1007 1 writedata5
rlabel metal2 2452 1008 2452 1008 1 writedata4
rlabel metal2 2152 1007 2152 1007 1 writedata3
rlabel metal2 1252 1006 1252 1006 1 writedata0
rlabel metal3 1006 3661 1006 3661 1 ph1
rlabel metal2 1006 3961 1006 3961 1 ph2
rlabel metal2 1261 3996 1261 3996 1 reset
rlabel metal2 1348 3996 1348 3996 1 adr0
rlabel metal2 1648 3996 1648 3996 1 adr1
rlabel metal2 1948 3995 1948 3995 1 adr2
rlabel metal2 2248 3995 2248 3995 1 adr3
rlabel metal2 2548 3995 2548 3995 1 adr4
rlabel metal2 2848 3996 2848 3996 1 adr5
rlabel metal2 3149 3996 3149 3996 1 adr6
rlabel metal2 3448 3996 3448 3996 1 adr7
rlabel metal2 3748 3996 3748 3996 1 memwrite
rlabel metal1 3995 3847 3995 3847 1 Vdd!
rlabel metal2 3994 3548 3994 3548 1 Gnd!
rlabel metal3 1004 1048 1004 1048 1 memdata0
rlabel metal3 1004 1348 1004 1348 1 memdata1
rlabel metal3 1005 1861 1005 1861 1 memdata2
rlabel metal3 1004 2161 1004 2161 1 memdata3
rlabel metal3 1004 2461 1004 2461 1 memdata4
rlabel metal3 1005 2761 1005 2761 1 memdata5
rlabel metal3 1005 3061 1005 3061 1 memdata6
rlabel metal3 1005 3361 1005 3361 1 memdata7
rlabel metal3 1972 2530 1972 2530 1 instr7
rlabel metal3 1973 2420 1973 2420 1 instr6
rlabel metal3 1973 2309 1973 2309 1 instr5
rlabel metal3 1973 2199 1973 2199 1 instr4
rlabel metal3 1973 2089 1973 2089 1 instr3
rlabel metal3 1973 1980 1973 1980 1 instr2
rlabel metal3 1973 1869 1973 1869 1 instr1
rlabel metal3 1974 1760 1974 1760 1 instr0
rlabel metal2 1449 1004 1449 1004 1 writedata1
rlabel metal2 1850 1005 1852 1007 1 writedata2
rlabel metal2 1698 3114 1698 3114 1 iord
rlabel metal1 1286 2516 1286 2516 1 pc7
rlabel metal3 1261 2508 1261 2508 1 aluout7
rlabel metal3 1261 2398 1261 2398 1 aluout6
rlabel metal1 1286 2406 1286 2406 1 pc6
rlabel metal3 1261 2289 1261 2289 1 aluout5
rlabel metal1 1286 2296 1286 2296 1 pc5
rlabel metal1 1286 2186 1286 2186 1 pc4
rlabel metal3 1261 2178 1261 2178 1 aluout4
rlabel metal1 1286 2075 1286 2075 1 pc3
rlabel metal3 1261 2068 1261 2068 1 aluout3
rlabel metal1 1286 1966 1286 1966 1 pc2
rlabel metal3 1261 1959 1261 1959 1 aluout2
rlabel metal1 1286 1856 1286 1856 1 pc1
rlabel metal3 1261 1849 1261 1849 1 aluout1
rlabel metal1 1286 1746 1286 1746 1 pc0
rlabel metal3 1261 1739 1261 1739 1 aluout0
rlabel metal2 3305 2571 3305 2571 1 pcen
rlabel metal1 3301 2514 3301 2514 1 pcnext7
rlabel metal1 3301 2404 3301 2404 1 pcnext6
rlabel metal1 3301 2294 3301 2294 1 pcnext5
rlabel metal1 3301 2184 3301 2184 1 pcnext4
rlabel metal1 3301 2074 3301 2074 1 pcnext3
rlabel metal1 3301 1964 3301 1964 1 pcnext2
rlabel metal1 3301 1854 3301 1854 1 pcnext1
rlabel metal1 3299 1744 3299 1744 1 pcnext0
rlabel metal2 3249 3006 3249 3006 1 pcsrc1
rlabel metal2 3217 3006 3217 3006 1 pcsrc0
rlabel metal3 3826 2508 3826 2508 1 aluresult7
rlabel metal3 3817 2397 3817 2397 1 aluresult6
rlabel metal3 3814 2277 3814 2277 1 aluresult5
rlabel metal3 3814 2167 3814 2167 1 aluresult4
rlabel metal3 3817 2050 3817 2050 1 aluresult3
rlabel metal3 3815 1957 3815 1957 1 aluresult2
rlabel metal3 3817 1836 3817 1836 1 aluresult1
rlabel metal3 3813 1738 3813 1738 1 aluresult0
<< end >>
