magic
tech scmos
timestamp 1493138306
<< m2contact >>
rect 6 12 10 16
<< metal2 >>
rect 22 64 26 65
rect 6 32 10 47
rect 14 41 18 46
rect 22 42 26 60
rect 30 42 34 46
rect 14 36 18 37
rect 54 0 58 112
rect 62 0 66 112
rect 70 32 74 57
rect 70 27 74 28
rect 94 0 98 112
rect 110 0 114 112
rect 182 106 186 112
rect 174 102 186 106
rect 158 65 162 66
rect 158 59 162 61
rect 174 65 178 102
rect 158 51 162 52
rect 134 47 138 48
rect 134 41 138 43
rect 142 32 146 40
rect 142 27 146 28
rect 174 2 178 61
rect 182 56 186 98
rect 270 65 274 112
rect 182 0 186 52
rect 230 7 234 61
rect 294 56 298 112
rect 310 87 314 112
rect 237 38 241 43
rect 270 29 274 52
rect 286 47 290 56
rect 286 38 290 43
rect 230 2 234 3
rect 270 7 274 9
rect 270 0 274 3
rect 294 0 298 25
rect 302 6 306 83
rect 310 82 314 83
rect 310 6 314 8
rect 310 0 314 2
rect 318 0 322 112
rect 350 60 354 61
rect 326 16 330 56
<< m3contact >>
rect 6 60 10 64
rect 22 60 26 64
rect 6 47 10 51
rect 30 46 34 50
rect 38 46 42 50
rect 14 37 18 41
rect 6 28 10 32
rect 6 12 10 16
rect 86 38 90 42
rect 70 28 74 32
rect 118 60 122 64
rect 158 61 162 65
rect 174 61 178 65
rect 158 52 162 56
rect 134 43 138 47
rect 150 43 154 47
rect 142 28 146 32
rect 182 52 186 56
rect 230 61 234 65
rect 270 61 274 65
rect 270 52 274 56
rect 237 43 241 47
rect 246 43 250 47
rect 237 34 241 38
rect 294 52 298 56
rect 302 83 306 87
rect 286 43 290 47
rect 270 25 274 29
rect 294 25 298 29
rect 230 3 234 7
rect 270 3 274 7
rect 310 83 314 87
rect 302 2 306 6
rect 310 2 314 6
rect 350 61 354 65
rect 366 41 370 45
rect 326 12 330 16
<< metal3 >>
rect 301 87 315 88
rect 301 83 302 87
rect 306 83 310 87
rect 314 83 315 87
rect 301 82 315 83
rect 157 65 179 66
rect 5 64 123 65
rect 5 60 6 64
rect 10 60 22 64
rect 26 60 118 64
rect 122 60 123 64
rect 157 61 158 65
rect 162 61 174 65
rect 178 61 179 65
rect 157 60 179 61
rect 229 65 355 66
rect 229 61 230 65
rect 234 61 270 65
rect 274 61 350 65
rect 354 61 355 65
rect 229 60 355 61
rect 5 59 123 60
rect 157 56 187 57
rect 157 52 158 56
rect 162 52 182 56
rect 186 52 187 56
rect 5 51 11 52
rect 157 51 187 52
rect 269 56 299 57
rect 269 52 270 56
rect 274 52 294 56
rect 298 52 299 56
rect 269 51 299 52
rect 5 47 6 51
rect 10 47 11 51
rect 5 46 11 47
rect 29 50 43 51
rect 29 46 30 50
rect 34 46 38 50
rect 42 46 43 50
rect 29 45 43 46
rect 133 47 242 48
rect 133 43 134 47
rect 138 43 150 47
rect 154 43 237 47
rect 241 43 242 47
rect 85 42 91 43
rect 133 42 242 43
rect 245 47 291 48
rect 245 43 246 47
rect 250 43 286 47
rect 290 43 291 47
rect 245 42 291 43
rect 365 45 371 46
rect 13 41 86 42
rect 13 37 14 41
rect 18 38 86 41
rect 90 38 91 42
rect 365 41 366 45
rect 370 41 371 45
rect 365 40 371 41
rect 18 37 91 38
rect 13 36 91 37
rect 236 38 299 39
rect 236 34 237 38
rect 241 34 299 38
rect 236 33 299 34
rect 5 32 147 33
rect 5 28 6 32
rect 10 28 70 32
rect 74 28 142 32
rect 146 28 147 32
rect 5 27 147 28
rect 269 29 299 30
rect 269 25 270 29
rect 274 25 294 29
rect 298 25 299 29
rect 269 24 299 25
rect 5 16 331 17
rect 5 12 6 16
rect 10 12 326 16
rect 330 12 331 16
rect 5 11 331 12
rect 229 7 275 8
rect 229 3 230 7
rect 234 3 270 7
rect 274 3 275 7
rect 229 2 275 3
rect 301 6 315 7
rect 301 2 302 6
rect 306 2 310 6
rect 314 2 315 6
rect 301 1 315 2
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 6 0 1 4
box -6 -4 18 96
use inv_1x  inv_1x_1
timestamp 1484418501
transform 1 0 22 0 1 4
box -6 -4 18 96
use mux4_dp_1x  mux4_dp_1x_0
timestamp 1484419186
transform 1 0 38 0 1 4
box -6 -4 106 96
use fulladder  fulladder_0
timestamp 1484419411
transform 1 0 144 0 1 4
box -8 -4 128 96
use mux4_dp_1x  mux4_dp_1x_1
timestamp 1484419186
transform 1 0 270 0 1 4
box -6 -4 106 96
<< labels >>
rlabel m3contact 8 62 8 62 1 B
rlabel m3contact 8 49 8 49 1 A
rlabel m3contact 8 14 8 14 1 Less
rlabel metal2 56 110 56 110 5 op6
rlabel metal2 64 110 64 110 5 op5
rlabel metal2 96 110 96 110 5 op4
rlabel metal2 112 110 112 110 5 op3
rlabel metal2 272 110 272 110 5 op0
rlabel metal2 296 110 296 110 5 op0b
rlabel metal2 312 110 312 110 5 op1
rlabel metal2 320 110 320 110 5 op1b
rlabel m3contact 248 45 248 45 1 y_temp
rlabel metal2 184 109 184 109 5 cout
rlabel metal3 368 46 368 46 1 result
<< end >>
