magic
tech scmos
timestamp 1492530230
<< metal1 >>
rect 30 325 666 340
rect 55 300 641 315
rect 55 287 641 293
rect 178 248 182 257
rect 490 251 493 256
rect 474 248 493 251
rect 314 233 318 242
rect 482 240 501 243
rect 138 198 150 202
rect 30 187 666 193
rect 338 128 373 131
rect 307 125 317 128
rect 386 123 390 132
rect 55 87 641 93
rect 55 65 641 80
rect 30 40 666 55
<< metal2 >>
rect 30 40 45 340
rect 55 65 70 315
rect 82 251 85 321
rect 98 228 101 301
rect 90 198 101 201
rect 98 141 101 198
rect 98 138 109 141
rect 106 125 109 138
rect 114 135 117 211
rect 122 178 125 231
rect 130 130 133 251
rect 154 228 157 244
rect 162 208 165 254
rect 178 248 181 271
rect 186 198 189 241
rect 194 198 197 231
rect 218 228 221 281
rect 234 251 237 261
rect 258 253 261 271
rect 298 251 301 271
rect 226 198 229 211
rect 242 198 245 231
rect 138 118 141 131
rect 202 121 205 141
rect 210 135 213 191
rect 266 178 269 201
rect 306 198 309 241
rect 314 238 349 241
rect 322 221 325 231
rect 314 218 325 221
rect 290 148 293 181
rect 226 108 229 132
rect 234 118 237 131
rect 314 125 317 218
rect 330 198 333 231
rect 338 168 341 221
rect 346 188 349 238
rect 370 138 373 251
rect 394 228 397 244
rect 370 135 381 138
rect 338 118 341 131
rect 394 129 397 141
rect 402 125 405 254
rect 426 251 429 261
rect 434 257 437 271
rect 474 231 477 251
rect 466 228 477 231
rect 418 188 421 201
rect 466 125 469 228
rect 482 201 485 241
rect 490 221 493 241
rect 490 218 501 221
rect 522 218 525 251
rect 578 228 581 251
rect 482 198 493 201
rect 490 137 493 198
rect 474 108 477 132
rect 498 128 501 218
rect 490 88 493 111
rect 506 58 509 201
rect 554 118 557 131
rect 562 129 565 151
rect 570 111 573 201
rect 586 188 589 231
rect 578 111 581 132
rect 586 123 589 141
rect 562 98 565 111
rect 570 108 581 111
rect 626 65 641 315
rect 651 40 666 340
<< metal3 >>
rect 0 317 86 322
rect 0 297 102 302
rect 0 277 302 282
rect 297 272 302 277
rect 97 267 262 272
rect 297 267 438 272
rect 0 257 566 262
rect 81 247 342 252
rect 441 247 606 252
rect 137 237 494 242
rect 513 237 574 242
rect 0 227 126 232
rect 153 227 470 232
rect 265 217 318 222
rect 337 217 390 222
rect 497 217 526 222
rect 113 207 374 212
rect 401 207 598 212
rect 0 197 142 202
rect 193 197 270 202
rect 305 197 494 202
rect 305 192 310 197
rect 209 187 310 192
rect 345 187 590 192
rect 265 177 294 182
rect 0 167 342 172
rect 129 157 406 162
rect 0 147 222 152
rect 489 147 566 152
rect 105 137 590 142
rect 0 127 390 132
rect 137 117 558 122
rect 225 107 574 112
rect 0 97 566 102
rect 417 87 494 92
rect 417 82 422 87
rect 0 77 422 82
rect 0 57 510 62
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1492530230
transform 1 0 37 0 1 332
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1492530230
transform 1 0 658 0 1 332
box -7 -7 7 7
use $$M3_M2  $$M3_M2_0
timestamp 1492530230
transform 1 0 84 0 1 320
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1492530230
transform 1 0 62 0 1 307
box -7 -7 7 7
use $$M3_M2  $$M3_M2_1
timestamp 1492530230
transform 1 0 100 0 1 300
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1492530230
transform 1 0 633 0 1 307
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1492530230
transform 1 0 62 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_2
timestamp 1492530230
transform 1 0 100 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1492530230
transform 1 0 84 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1492530230
transform 1 0 84 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_1
timestamp 1492530230
transform 1 0 100 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_6
timestamp 1492530230
transform 1 0 92 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_3
timestamp 1492530230
transform 1 0 132 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_5
timestamp 1492530230
transform 1 0 124 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_7
timestamp 1492530230
transform 1 0 116 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1492530230
transform 1 0 164 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_4
timestamp 1492530230
transform 1 0 140 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_5
timestamp 1492530230
transform 1 0 156 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1492530230
transform 1 0 140 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_6
timestamp 1492530230
transform 1 0 156 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_8
timestamp 1492530230
transform 1 0 164 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_7
timestamp 1492530230
transform 1 0 140 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1492530230
transform 1 0 140 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_11
timestamp 1492530230
transform 1 0 180 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_8
timestamp 1492530230
transform 1 0 180 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_12
timestamp 1492530230
transform 1 0 188 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_10
timestamp 1492530230
transform 1 0 196 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1492530230
transform 1 0 188 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1492530230
transform 1 0 196 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_10
timestamp 1492530230
transform 1 0 220 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1492530230
transform 1 0 220 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_13
timestamp 1492530230
transform 1 0 236 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_9
timestamp 1492530230
transform 1 0 236 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_12
timestamp 1492530230
transform 1 0 244 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_14
timestamp 1492530230
transform 1 0 228 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_14
timestamp 1492530230
transform 1 0 228 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_16
timestamp 1492530230
transform 1 0 244 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_18
timestamp 1492530230
transform 1 0 260 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_15
timestamp 1492530230
transform 1 0 260 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_16
timestamp 1492530230
transform 1 0 252 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_19
timestamp 1492530230
transform 1 0 252 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_17
timestamp 1492530230
transform 1 0 268 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_20
timestamp 1492530230
transform 1 0 268 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1492530230
transform 1 0 268 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_22
timestamp 1492530230
transform 1 0 300 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_18
timestamp 1492530230
transform 1 0 300 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_20
timestamp 1492530230
transform 1 0 308 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_21
timestamp 1492530230
transform 1 0 316 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_19
timestamp 1492530230
transform 1 0 340 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_23
timestamp 1492530230
transform 1 0 340 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_22
timestamp 1492530230
transform 1 0 324 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_24
timestamp 1492530230
transform 1 0 332 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_25
timestamp 1492530230
transform 1 0 316 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_27
timestamp 1492530230
transform 1 0 308 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_26
timestamp 1492530230
transform 1 0 340 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_23
timestamp 1492530230
transform 1 0 332 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_25
timestamp 1492530230
transform 1 0 372 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_24
timestamp 1492530230
transform 1 0 404 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_27
timestamp 1492530230
transform 1 0 380 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_26
timestamp 1492530230
transform 1 0 396 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_29
timestamp 1492530230
transform 1 0 380 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_30
timestamp 1492530230
transform 1 0 396 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_28
timestamp 1492530230
transform 1 0 388 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_31
timestamp 1492530230
transform 1 0 388 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_32
timestamp 1492530230
transform 1 0 372 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_33
timestamp 1492530230
transform 1 0 404 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_31
timestamp 1492530230
transform 1 0 420 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_34
timestamp 1492530230
transform 1 0 436 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_35
timestamp 1492530230
transform 1 0 428 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_29
timestamp 1492530230
transform 1 0 436 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_30
timestamp 1492530230
transform 1 0 428 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_32
timestamp 1492530230
transform 1 0 444 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_37
timestamp 1492530230
transform 1 0 444 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_33
timestamp 1492530230
transform 1 0 476 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_40
timestamp 1492530230
transform 1 0 468 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_34
timestamp 1492530230
transform 1 0 524 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_36
timestamp 1492530230
transform 1 0 484 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_38
timestamp 1492530230
transform 1 0 492 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_35
timestamp 1492530230
transform 1 0 516 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_39
timestamp 1492530230
transform 1 0 516 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_41
timestamp 1492530230
transform 1 0 500 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_42
timestamp 1492530230
transform 1 0 524 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_43
timestamp 1492530230
transform 1 0 492 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1492530230
transform 1 0 508 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_38
timestamp 1492530230
transform 1 0 564 0 1 259
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1492530230
transform 1 0 564 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_45
timestamp 1492530230
transform 1 0 580 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_40
timestamp 1492530230
transform 1 0 572 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_47
timestamp 1492530230
transform 1 0 572 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_41
timestamp 1492530230
transform 1 0 580 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_42
timestamp 1492530230
transform 1 0 588 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_43
timestamp 1492530230
transform 1 0 572 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1492530230
transform 1 0 604 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_46
timestamp 1492530230
transform 1 0 604 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1492530230
transform 1 0 596 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1492530230
transform 1 0 596 0 1 210
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1492530230
transform 1 0 633 0 1 290
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1492530230
transform 1 0 37 0 1 190
box -7 -2 7 2
use NAND2X1  NAND2X1_0
timestamp 1492530230
transform 1 0 80 0 -1 290
box -8 -3 32 105
use FILL  FILL_0
timestamp 1492530230
transform 1 0 104 0 -1 290
box -8 -3 16 105
use FILL  FILL_1
timestamp 1492530230
transform 1 0 112 0 -1 290
box -8 -3 16 105
use FILL  FILL_2
timestamp 1492530230
transform 1 0 120 0 -1 290
box -8 -3 16 105
use OAI22X1  OAI22X1_0
timestamp 1492530230
transform -1 0 168 0 -1 290
box -8 -3 46 105
use FILL  FILL_3
timestamp 1492530230
transform 1 0 168 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1492530230
transform 1 0 176 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_17
timestamp 1492530230
transform 1 0 212 0 1 190
box -3 -3 3 3
use FILL  FILL_4
timestamp 1492530230
transform 1 0 200 0 -1 290
box -8 -3 16 105
use FILL  FILL_5
timestamp 1492530230
transform 1 0 208 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1492530230
transform -1 0 240 0 -1 290
box -8 -3 32 105
use INVX2  INVX2_0
timestamp 1492530230
transform -1 0 256 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1492530230
transform 1 0 256 0 -1 290
box -9 -3 26 105
use FILL  FILL_6
timestamp 1492530230
transform 1 0 272 0 -1 290
box -8 -3 16 105
use FILL  FILL_7
timestamp 1492530230
transform 1 0 280 0 -1 290
box -8 -3 16 105
use FILL  FILL_8
timestamp 1492530230
transform 1 0 288 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1492530230
transform 1 0 296 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_28
timestamp 1492530230
transform 1 0 348 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_4
timestamp 1492530230
transform -1 0 344 0 -1 290
box -8 -3 32 105
use FILL  FILL_9
timestamp 1492530230
transform 1 0 344 0 -1 290
box -8 -3 16 105
use FILL  FILL_10
timestamp 1492530230
transform 1 0 352 0 -1 290
box -8 -3 16 105
use FILL  FILL_11
timestamp 1492530230
transform 1 0 360 0 -1 290
box -8 -3 16 105
use OAI22X1  OAI22X1_1
timestamp 1492530230
transform -1 0 408 0 -1 290
box -8 -3 46 105
use $$M3_M2  $$M3_M2_36
timestamp 1492530230
transform 1 0 420 0 1 190
box -3 -3 3 3
use FILL  FILL_12
timestamp 1492530230
transform 1 0 408 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1492530230
transform -1 0 432 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1492530230
transform 1 0 432 0 -1 290
box -9 -3 26 105
use FILL  FILL_13
timestamp 1492530230
transform 1 0 448 0 -1 290
box -8 -3 16 105
use FILL  FILL_14
timestamp 1492530230
transform 1 0 456 0 -1 290
box -8 -3 16 105
use FILL  FILL_15
timestamp 1492530230
transform 1 0 464 0 -1 290
box -8 -3 16 105
use FILL  FILL_16
timestamp 1492530230
transform 1 0 472 0 -1 290
box -8 -3 16 105
use FILL  FILL_17
timestamp 1492530230
transform 1 0 480 0 -1 290
box -8 -3 16 105
use OAI22X1  OAI22X1_2
timestamp 1492530230
transform 1 0 488 0 -1 290
box -8 -3 46 105
use FILL  FILL_18
timestamp 1492530230
transform 1 0 528 0 -1 290
box -8 -3 16 105
use FILL  FILL_19
timestamp 1492530230
transform 1 0 536 0 -1 290
box -8 -3 16 105
use FILL  FILL_20
timestamp 1492530230
transform 1 0 544 0 -1 290
box -8 -3 16 105
use FILL  FILL_21
timestamp 1492530230
transform 1 0 552 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_49
timestamp 1492530230
transform 1 0 588 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_5
timestamp 1492530230
transform 1 0 560 0 -1 290
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1492530230
transform -1 0 608 0 -1 290
box -8 -3 32 105
use FILL  FILL_22
timestamp 1492530230
transform 1 0 608 0 -1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1492530230
transform 1 0 658 0 1 190
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1492530230
transform 1 0 62 0 1 90
box -7 -2 7 2
use FILL  FILL_23
timestamp 1492530230
transform -1 0 88 0 1 90
box -8 -3 16 105
use FILL  FILL_24
timestamp 1492530230
transform -1 0 96 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_45
timestamp 1492530230
transform 1 0 124 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_50
timestamp 1492530230
transform 1 0 132 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_51
timestamp 1492530230
transform 1 0 108 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_46
timestamp 1492530230
transform 1 0 116 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_47
timestamp 1492530230
transform 1 0 132 0 1 132
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1492530230
transform 1 0 108 0 1 127
box -2 -2 2 2
use FILL  FILL_25
timestamp 1492530230
transform -1 0 104 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_48
timestamp 1492530230
transform 1 0 140 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_52
timestamp 1492530230
transform 1 0 140 0 1 120
box -3 -3 3 3
use OAI22X1  OAI22X1_3
timestamp 1492530230
transform 1 0 104 0 1 90
box -8 -3 46 105
use FILL  FILL_26
timestamp 1492530230
transform -1 0 152 0 1 90
box -8 -3 16 105
use FILL  FILL_27
timestamp 1492530230
transform -1 0 160 0 1 90
box -8 -3 16 105
use FILL  FILL_28
timestamp 1492530230
transform -1 0 168 0 1 90
box -8 -3 16 105
use FILL  FILL_29
timestamp 1492530230
transform -1 0 176 0 1 90
box -8 -3 16 105
use FILL  FILL_30
timestamp 1492530230
transform -1 0 184 0 1 90
box -8 -3 16 105
use FILL  FILL_31
timestamp 1492530230
transform -1 0 192 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_50
timestamp 1492530230
transform 1 0 220 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_55
timestamp 1492530230
transform 1 0 220 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_56
timestamp 1492530230
transform 1 0 204 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_51
timestamp 1492530230
transform 1 0 212 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_52
timestamp 1492530230
transform 1 0 228 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_54
timestamp 1492530230
transform 1 0 204 0 1 123
box -2 -2 2 2
use FILL  FILL_32
timestamp 1492530230
transform -1 0 200 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_53
timestamp 1492530230
transform 1 0 236 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_57
timestamp 1492530230
transform 1 0 236 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_58
timestamp 1492530230
transform 1 0 228 0 1 110
box -3 -3 3 3
use OAI22X1  OAI22X1_4
timestamp 1492530230
transform 1 0 200 0 1 90
box -8 -3 46 105
use FILL  FILL_33
timestamp 1492530230
transform -1 0 248 0 1 90
box -8 -3 16 105
use FILL  FILL_34
timestamp 1492530230
transform -1 0 256 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_53
timestamp 1492530230
transform 1 0 268 0 1 180
box -3 -3 3 3
use FILL  FILL_35
timestamp 1492530230
transform -1 0 264 0 1 90
box -8 -3 16 105
use FILL  FILL_36
timestamp 1492530230
transform -1 0 272 0 1 90
box -8 -3 16 105
use FILL  FILL_37
timestamp 1492530230
transform -1 0 280 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_54
timestamp 1492530230
transform 1 0 292 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_55
timestamp 1492530230
transform 1 0 292 0 1 150
box -2 -2 2 2
use FILL  FILL_38
timestamp 1492530230
transform -1 0 288 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_62
timestamp 1492530230
transform 1 0 300 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1492530230
transform 1 0 300 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_60
timestamp 1492530230
transform 1 0 316 0 1 127
box -2 -2 2 2
use NAND2X1  NAND2X1_7
timestamp 1492530230
transform -1 0 312 0 1 90
box -8 -3 32 105
use FILL  FILL_39
timestamp 1492530230
transform -1 0 320 0 1 90
box -8 -3 16 105
use FILL  FILL_40
timestamp 1492530230
transform -1 0 328 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_59
timestamp 1492530230
transform 1 0 340 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_58
timestamp 1492530230
transform 1 0 340 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_64
timestamp 1492530230
transform 1 0 340 0 1 120
box -3 -3 3 3
use FILL  FILL_41
timestamp 1492530230
transform -1 0 336 0 1 90
box -8 -3 16 105
use FILL  FILL_42
timestamp 1492530230
transform -1 0 344 0 1 90
box -8 -3 16 105
use FILL  FILL_43
timestamp 1492530230
transform -1 0 352 0 1 90
box -8 -3 16 105
use FILL  FILL_44
timestamp 1492530230
transform -1 0 360 0 1 90
box -8 -3 16 105
use FILL  FILL_45
timestamp 1492530230
transform -1 0 368 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_60
timestamp 1492530230
transform 1 0 404 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_56
timestamp 1492530230
transform 1 0 380 0 1 137
box -2 -2 2 2
use $$M3_M2  $$M3_M2_61
timestamp 1492530230
transform 1 0 396 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1492530230
transform 1 0 388 0 1 130
box -2 -2 2 2
use $$M2_M1  $$M2_M1_57
timestamp 1492530230
transform 1 0 396 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1492530230
transform 1 0 388 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1492530230
transform 1 0 404 0 1 127
box -2 -2 2 2
use OAI22X1  OAI22X1_5
timestamp 1492530230
transform -1 0 408 0 1 90
box -8 -3 46 105
use FILL  FILL_46
timestamp 1492530230
transform -1 0 416 0 1 90
box -8 -3 16 105
use FILL  FILL_47
timestamp 1492530230
transform -1 0 424 0 1 90
box -8 -3 16 105
use FILL  FILL_48
timestamp 1492530230
transform -1 0 432 0 1 90
box -8 -3 16 105
use FILL  FILL_49
timestamp 1492530230
transform -1 0 440 0 1 90
box -8 -3 16 105
use FILL  FILL_50
timestamp 1492530230
transform -1 0 448 0 1 90
box -8 -3 16 105
use FILL  FILL_51
timestamp 1492530230
transform -1 0 456 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_65
timestamp 1492530230
transform 1 0 492 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_63
timestamp 1492530230
transform 1 0 492 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_64
timestamp 1492530230
transform 1 0 476 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_66
timestamp 1492530230
transform 1 0 468 0 1 127
box -2 -2 2 2
use FILL  FILL_52
timestamp 1492530230
transform -1 0 464 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_65
timestamp 1492530230
transform 1 0 500 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_66
timestamp 1492530230
transform 1 0 476 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_67
timestamp 1492530230
transform 1 0 492 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1492530230
transform 1 0 492 0 1 90
box -3 -3 3 3
use OAI22X1  OAI22X1_6
timestamp 1492530230
transform 1 0 464 0 1 90
box -8 -3 46 105
use FILL  FILL_53
timestamp 1492530230
transform -1 0 512 0 1 90
box -8 -3 16 105
use FILL  FILL_54
timestamp 1492530230
transform -1 0 520 0 1 90
box -8 -3 16 105
use FILL  FILL_55
timestamp 1492530230
transform -1 0 528 0 1 90
box -8 -3 16 105
use FILL  FILL_56
timestamp 1492530230
transform -1 0 536 0 1 90
box -8 -3 16 105
use FILL  FILL_57
timestamp 1492530230
transform -1 0 544 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_67
timestamp 1492530230
transform 1 0 564 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_68
timestamp 1492530230
transform 1 0 588 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_70
timestamp 1492530230
transform 1 0 556 0 1 130
box -2 -2 2 2
use $$M2_M1  $$M2_M1_68
timestamp 1492530230
transform 1 0 564 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_69
timestamp 1492530230
transform 1 0 580 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_69
timestamp 1492530230
transform 1 0 556 0 1 120
box -3 -3 3 3
use FILL  FILL_58
timestamp 1492530230
transform -1 0 552 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_71
timestamp 1492530230
transform 1 0 588 0 1 124
box -2 -2 2 2
use $$M2_M1  $$M2_M1_72
timestamp 1492530230
transform 1 0 564 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_70
timestamp 1492530230
transform 1 0 572 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_71
timestamp 1492530230
transform 1 0 564 0 1 100
box -3 -3 3 3
use OAI22X1  OAI22X1_7
timestamp 1492530230
transform -1 0 592 0 1 90
box -8 -3 46 105
use FILL  FILL_59
timestamp 1492530230
transform -1 0 600 0 1 90
box -8 -3 16 105
use FILL  FILL_60
timestamp 1492530230
transform -1 0 608 0 1 90
box -8 -3 16 105
use FILL  FILL_61
timestamp 1492530230
transform -1 0 616 0 1 90
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1492530230
transform 1 0 633 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1492530230
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1492530230
transform 1 0 633 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_73
timestamp 1492530230
transform 1 0 508 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1492530230
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1492530230
transform 1 0 658 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 260 2 260 4 FreeSans 26 0 0 0 right
flabel metal3 2 280 2 280 4 FreeSans 26 0 0 0 k[2]
flabel metal3 2 320 2 320 4 FreeSans 26 0 0 0 k[1]
flabel metal3 2 300 2 300 4 FreeSans 26 0 0 0 k[0]
flabel metal3 2 150 2 150 4 FreeSans 26 0 0 0 s[0]
flabel metal3 2 80 2 80 4 FreeSans 26 0 0 0 s[2]
flabel metal3 2 100 2 100 4 FreeSans 26 0 0 0 s[3]
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 s[1]
flabel metal3 2 230 2 230 4 FreeSans 26 0 0 0 s[7]
flabel metal3 2 130 2 130 4 FreeSans 26 0 0 0 s[4]
flabel metal3 2 170 2 170 4 FreeSans 26 0 0 0 s[5]
flabel metal3 2 200 2 200 4 FreeSans 26 0 0 0 s[6]
rlabel metal1 170 334 170 334 1 Vdd!
rlabel metal1 169 308 169 308 1 Gnd!
<< end >>
