magic
tech scmos
timestamp 1492530230
<< m2contact >>
rect -7 -2 7 2
<< end >>
