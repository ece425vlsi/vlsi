magic
tech scmos
timestamp 1493747787
<< metal2 >>
rect 1670 1953 1826 1957
rect 564 1941 568 1942
rect 380 1932 384 1933
rect 364 1923 368 1924
rect 356 1914 360 1915
rect 348 1905 352 1906
rect 340 1896 344 1897
rect 332 1887 336 1888
rect 324 1878 328 1879
rect 196 1869 200 1870
rect 140 1860 144 1861
rect 196 1859 200 1865
rect 324 1856 328 1874
rect 332 1858 336 1883
rect 340 1856 344 1892
rect 348 1856 352 1901
rect 356 1855 360 1910
rect 364 1856 368 1919
rect 380 1853 384 1928
rect 564 1854 568 1937
rect 581 1860 585 1952
rect 605 1869 609 1952
rect 637 1878 641 1952
rect 669 1887 673 1952
rect 709 1896 713 1952
rect 741 1905 745 1952
rect 773 1914 777 1952
rect 805 1923 809 1952
rect 837 1932 841 1952
rect 869 1941 873 1952
rect 869 1936 873 1937
rect 837 1927 841 1928
rect 852 1932 856 1933
rect 805 1918 809 1919
rect 836 1923 840 1924
rect 773 1909 777 1910
rect 741 1900 745 1901
rect 709 1891 713 1892
rect 724 1896 728 1897
rect 669 1882 673 1883
rect 637 1873 641 1874
rect 605 1864 609 1865
rect 724 1859 728 1892
rect 836 1856 840 1919
rect 852 1858 856 1928
rect 860 1914 864 1915
rect 860 1859 864 1910
rect 868 1905 872 1906
rect 868 1856 872 1901
rect 909 1896 913 1952
rect 941 1923 945 1952
rect 973 1932 977 1952
rect 973 1927 977 1928
rect 941 1918 945 1919
rect 1005 1914 1009 1952
rect 1005 1909 1009 1910
rect 1037 1905 1041 1952
rect 1037 1900 1041 1901
rect 909 1891 913 1892
rect 932 1896 936 1897
rect 876 1887 880 1888
rect 876 1859 880 1883
rect 884 1878 888 1879
rect 884 1859 888 1874
rect 892 1869 896 1870
rect 892 1859 896 1865
rect 932 1859 936 1892
rect 1069 1887 1073 1952
rect 1069 1882 1073 1883
rect 1109 1878 1113 1952
rect 1109 1873 1113 1874
rect 1141 1869 1145 1952
rect 1173 1896 1177 1952
rect 1173 1891 1177 1892
rect 1141 1864 1145 1865
rect 1100 1860 1104 1861
rect 1100 1854 1104 1856
rect 1205 1860 1209 1952
rect 1205 1855 1209 1856
rect 1237 1860 1241 1952
rect 1269 1869 1273 1952
rect 1309 1879 1313 1952
rect 1341 1888 1345 1952
rect 1373 1897 1377 1952
rect 1405 1906 1409 1952
rect 1437 1915 1441 1952
rect 1469 1924 1473 1952
rect 1509 1933 1513 1952
rect 1541 1942 1545 1952
rect 1573 1951 1577 1952
rect 1573 1946 1577 1947
rect 1606 1943 1609 1953
rect 1638 1950 1641 1952
rect 1638 1946 1818 1950
rect 1606 1939 1810 1943
rect 1541 1937 1545 1938
rect 1509 1928 1513 1929
rect 1469 1919 1473 1920
rect 1437 1910 1441 1911
rect 1405 1901 1409 1902
rect 1373 1892 1377 1893
rect 1341 1883 1345 1884
rect 1772 1888 1776 1889
rect 1309 1874 1313 1875
rect 1740 1879 1744 1880
rect 1269 1864 1273 1865
rect 1724 1869 1728 1870
rect 1237 1855 1241 1856
rect 1636 1860 1640 1861
rect 1724 1856 1728 1865
rect 1740 1856 1744 1875
rect 1772 1857 1776 1884
rect 1806 1860 1810 1939
rect 1814 1869 1818 1946
rect 1822 1878 1826 1953
rect 2421 1951 2425 1952
rect 2389 1942 2393 1943
rect 2381 1933 2385 1934
rect 2188 1924 2192 1925
rect 2132 1915 2136 1916
rect 2100 1906 2104 1907
rect 1822 1873 1826 1874
rect 1948 1897 1952 1898
rect 1814 1864 1818 1865
rect 1948 1860 1952 1893
rect 2100 1860 2104 1902
rect 2132 1860 2136 1911
rect 2188 1858 2192 1920
rect 2381 1860 2385 1929
rect 2389 1860 2393 1938
rect 2421 1859 2425 1947
rect 2733 1878 2737 1879
rect 2637 1869 2641 1870
rect 2637 1860 2641 1865
rect 2733 1861 2737 1874
rect 1636 1855 1640 1856
rect 1806 1855 1810 1856
<< m3contact >>
rect 564 1937 568 1941
rect 380 1928 384 1932
rect 364 1919 368 1923
rect 356 1910 360 1914
rect 348 1901 352 1905
rect 340 1892 344 1896
rect 332 1883 336 1887
rect 324 1874 328 1878
rect 196 1865 200 1869
rect 140 1856 144 1860
rect 869 1937 873 1941
rect 837 1928 841 1932
rect 852 1928 856 1932
rect 805 1919 809 1923
rect 836 1919 840 1923
rect 773 1910 777 1914
rect 741 1901 745 1905
rect 709 1892 713 1896
rect 724 1892 728 1896
rect 669 1883 673 1887
rect 637 1874 641 1878
rect 605 1865 609 1869
rect 581 1856 585 1860
rect 860 1910 864 1914
rect 868 1901 872 1905
rect 973 1928 977 1932
rect 941 1919 945 1923
rect 1005 1910 1009 1914
rect 1037 1901 1041 1905
rect 909 1892 913 1896
rect 932 1892 936 1896
rect 876 1883 880 1887
rect 884 1874 888 1878
rect 892 1865 896 1869
rect 1069 1883 1073 1887
rect 1109 1874 1113 1878
rect 1173 1892 1177 1896
rect 1141 1865 1145 1869
rect 1100 1856 1104 1860
rect 1205 1856 1209 1860
rect 1573 1947 1577 1951
rect 1541 1938 1545 1942
rect 1509 1929 1513 1933
rect 1469 1920 1473 1924
rect 1437 1911 1441 1915
rect 1405 1902 1409 1906
rect 1373 1893 1377 1897
rect 1341 1884 1345 1888
rect 1772 1884 1776 1888
rect 1309 1875 1313 1879
rect 1740 1875 1744 1879
rect 1269 1865 1273 1869
rect 1724 1865 1728 1869
rect 1237 1856 1241 1860
rect 1636 1856 1640 1860
rect 2421 1947 2425 1951
rect 2389 1938 2393 1942
rect 2381 1929 2385 1933
rect 2188 1920 2192 1924
rect 2132 1911 2136 1915
rect 2100 1902 2104 1906
rect 1822 1874 1826 1878
rect 1948 1893 1952 1897
rect 1814 1865 1818 1869
rect 1806 1856 1810 1860
rect 2733 1874 2737 1878
rect 2637 1865 2641 1869
rect 2597 1856 2601 1860
<< metal3 >>
rect 1572 1951 2426 1952
rect 1572 1947 1573 1951
rect 1577 1947 2421 1951
rect 2425 1947 2426 1951
rect 1572 1946 2426 1947
rect 1540 1942 2394 1943
rect 563 1941 874 1942
rect 563 1937 564 1941
rect 568 1937 869 1941
rect 873 1937 874 1941
rect 1540 1938 1541 1942
rect 1545 1938 2389 1942
rect 2393 1938 2394 1942
rect 1540 1937 2394 1938
rect 563 1936 874 1937
rect 1508 1933 2386 1934
rect 379 1932 842 1933
rect 379 1928 380 1932
rect 384 1928 837 1932
rect 841 1928 842 1932
rect 379 1927 842 1928
rect 851 1932 978 1933
rect 851 1928 852 1932
rect 856 1928 973 1932
rect 977 1928 978 1932
rect 1508 1929 1509 1933
rect 1513 1929 2381 1933
rect 2385 1929 2386 1933
rect 1508 1928 2386 1929
rect 851 1927 978 1928
rect 1468 1924 2193 1925
rect 363 1923 810 1924
rect 363 1919 364 1923
rect 368 1919 805 1923
rect 809 1919 810 1923
rect 363 1918 810 1919
rect 835 1923 946 1924
rect 835 1919 836 1923
rect 840 1919 941 1923
rect 945 1919 946 1923
rect 1468 1920 1469 1924
rect 1473 1920 2188 1924
rect 2192 1920 2193 1924
rect 1468 1919 2193 1920
rect 835 1918 946 1919
rect 1436 1915 2137 1916
rect 355 1914 778 1915
rect 355 1910 356 1914
rect 360 1910 773 1914
rect 777 1910 778 1914
rect 355 1909 778 1910
rect 859 1914 1010 1915
rect 859 1910 860 1914
rect 864 1910 1005 1914
rect 1009 1910 1010 1914
rect 1436 1911 1437 1915
rect 1441 1911 2132 1915
rect 2136 1911 2137 1915
rect 1436 1910 2137 1911
rect 859 1909 1010 1910
rect 1404 1906 2105 1907
rect 347 1905 746 1906
rect 347 1901 348 1905
rect 352 1901 741 1905
rect 745 1901 746 1905
rect 347 1900 746 1901
rect 867 1905 1042 1906
rect 867 1901 868 1905
rect 872 1901 1037 1905
rect 1041 1901 1042 1905
rect 1404 1902 1405 1906
rect 1409 1902 2100 1906
rect 2104 1902 2105 1906
rect 1404 1901 2105 1902
rect 867 1900 1042 1901
rect 1372 1897 1953 1898
rect 339 1896 714 1897
rect 339 1892 340 1896
rect 344 1892 709 1896
rect 713 1892 714 1896
rect 339 1891 714 1892
rect 723 1896 914 1897
rect 723 1892 724 1896
rect 728 1892 909 1896
rect 913 1892 914 1896
rect 723 1891 914 1892
rect 931 1896 1178 1897
rect 931 1892 932 1896
rect 936 1892 1173 1896
rect 1177 1892 1178 1896
rect 1372 1893 1373 1897
rect 1377 1893 1948 1897
rect 1952 1893 1953 1897
rect 1372 1892 1953 1893
rect 931 1891 1178 1892
rect 1340 1888 1777 1889
rect 331 1887 674 1888
rect 331 1883 332 1887
rect 336 1883 669 1887
rect 673 1883 674 1887
rect 331 1882 674 1883
rect 875 1887 1074 1888
rect 875 1883 876 1887
rect 880 1883 1069 1887
rect 1073 1883 1074 1887
rect 1340 1884 1341 1888
rect 1345 1884 1772 1888
rect 1776 1884 1777 1888
rect 1340 1883 1777 1884
rect 875 1882 1074 1883
rect 1308 1879 1745 1880
rect 323 1878 642 1879
rect 323 1874 324 1878
rect 328 1874 637 1878
rect 641 1874 642 1878
rect 323 1873 642 1874
rect 883 1878 1114 1879
rect 883 1874 884 1878
rect 888 1874 1109 1878
rect 1113 1874 1114 1878
rect 1308 1875 1309 1879
rect 1313 1875 1740 1879
rect 1744 1875 1745 1879
rect 1308 1874 1745 1875
rect 1821 1878 2738 1879
rect 1821 1874 1822 1878
rect 1826 1874 2733 1878
rect 2737 1874 2738 1878
rect 883 1873 1114 1874
rect 1821 1873 2738 1874
rect 195 1869 610 1870
rect 195 1865 196 1869
rect 200 1865 605 1869
rect 609 1865 610 1869
rect 195 1864 610 1865
rect 891 1869 1146 1870
rect 891 1865 892 1869
rect 896 1865 1141 1869
rect 1145 1865 1146 1869
rect 891 1864 1146 1865
rect 1268 1869 1729 1870
rect 1268 1865 1269 1869
rect 1273 1865 1724 1869
rect 1728 1865 1729 1869
rect 1268 1864 1729 1865
rect 1813 1869 2642 1870
rect 1813 1865 1814 1869
rect 1818 1865 2637 1869
rect 2641 1865 2642 1869
rect 1813 1864 2642 1865
rect 139 1860 586 1861
rect 139 1856 140 1860
rect 144 1856 581 1860
rect 585 1856 586 1860
rect 139 1855 586 1856
rect 1099 1860 1210 1861
rect 1099 1856 1100 1860
rect 1104 1856 1205 1860
rect 1209 1856 1210 1860
rect 1099 1855 1210 1856
rect 1236 1860 1641 1861
rect 1236 1856 1237 1860
rect 1241 1856 1636 1860
rect 1640 1856 1641 1860
rect 1236 1855 1641 1856
rect 1805 1860 2602 1861
rect 1805 1856 1806 1860
rect 1810 1856 2597 1860
rect 2601 1856 2602 1860
rect 1805 1855 2602 1856
use alt_controller  alt_controller_0
timestamp 1493747238
transform 1 0 540 0 1 1952
box 0 0 2082 380
use datapath  datapath_0
timestamp 1493747238
transform 1 0 140 0 1 548
box -140 -548 2736 1343
<< end >>
