magic
tech scmos
timestamp 1486491337
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 23
rect 10 7 12 23
rect 15 7 17 23
<< ptransistor >>
rect 5 70 7 83
rect 13 70 15 83
rect 21 70 23 83
<< ndiffusion >>
rect 0 22 5 23
rect 4 8 5 22
rect 0 7 5 8
rect 7 7 10 23
rect 12 7 15 23
rect 17 22 22 23
rect 17 8 18 22
rect 17 7 22 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 72 5 81
rect 0 70 5 72
rect 7 81 13 83
rect 7 72 8 81
rect 12 72 13 81
rect 7 70 13 72
rect 15 81 21 83
rect 15 72 16 81
rect 20 72 21 81
rect 15 70 21 72
rect 23 81 28 83
rect 23 72 24 81
rect 23 70 28 72
<< ndcontact >>
rect 0 8 4 22
rect 18 8 22 22
<< pdcontact >>
rect 0 72 4 81
rect 8 72 12 81
rect 16 72 20 81
rect 24 72 28 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 5 69 7 70
rect 13 69 15 70
rect 1 67 7 69
rect 10 67 15 69
rect 1 28 3 67
rect 1 26 7 28
rect 5 23 7 26
rect 10 23 12 67
rect 21 59 23 70
rect 20 57 23 59
rect 20 26 22 57
rect 15 24 22 26
rect 15 23 17 24
rect 5 5 7 7
rect 10 5 12 7
rect 15 5 17 7
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 81 4 86
rect 16 81 20 86
rect 0 70 4 72
rect 24 81 28 83
rect 8 66 12 72
rect 24 66 28 72
rect 8 62 28 66
rect 24 47 28 62
rect 24 23 28 43
rect 0 22 4 23
rect 0 4 4 8
rect 18 22 28 23
rect 22 19 28 22
rect 18 7 22 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
<< end >>
