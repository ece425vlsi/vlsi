magic
tech scmos
timestamp 1490995571
<< metal1 >>
rect 30 525 954 540
rect 55 500 929 515
rect 55 487 929 493
rect 98 478 117 481
rect 146 467 150 471
rect 146 464 157 467
rect 250 458 254 467
rect 315 461 325 464
rect 306 448 310 457
rect 346 453 350 462
rect 426 456 437 459
rect 683 458 693 461
rect 730 458 734 467
rect 618 451 629 454
rect 402 448 421 451
rect 482 447 493 450
rect 714 448 718 457
rect 117 428 121 436
rect 162 432 166 442
rect 402 438 413 441
rect 391 431 398 436
rect 410 435 413 438
rect 474 432 478 442
rect 707 438 725 441
rect 647 431 654 436
rect 802 434 806 442
rect 391 428 405 431
rect 507 428 517 431
rect 647 428 661 431
rect 258 398 267 402
rect 30 387 954 393
rect 450 358 454 368
rect 411 348 421 351
rect 578 348 589 351
rect 490 341 494 348
rect 655 344 662 352
rect 274 338 285 341
rect 490 338 501 341
rect 802 338 806 346
rect 202 330 229 333
rect 267 330 277 333
rect 458 331 469 334
rect 490 333 494 338
rect 498 334 501 338
rect 498 331 509 334
rect 386 327 397 330
rect 251 321 259 327
rect 314 321 341 324
rect 354 322 365 325
rect 530 323 534 332
rect 722 328 726 337
rect 195 318 205 321
rect 242 318 259 321
rect 402 313 411 321
rect 611 318 621 321
rect 55 287 929 293
rect 314 278 325 281
rect 105 257 110 261
rect 474 258 478 267
rect 342 255 357 258
rect 370 248 375 257
rect 514 248 518 257
rect 522 243 526 252
rect 561 248 566 257
rect 594 251 598 257
rect 578 248 598 251
rect 250 234 254 242
rect 362 228 369 236
rect 394 235 405 238
rect 482 232 486 242
rect 498 240 509 243
rect 602 242 621 245
rect 498 231 501 240
rect 627 238 637 241
rect 490 228 501 231
rect 567 228 574 236
rect 610 228 621 231
rect 674 228 681 236
rect 445 198 454 202
rect 30 187 954 193
rect 227 178 261 181
rect 587 178 597 181
rect 194 138 198 146
rect 426 133 430 142
rect 506 137 525 140
rect 530 138 534 148
rect 658 128 662 137
rect 778 128 901 131
rect 778 125 782 128
rect 410 119 415 123
rect 738 118 773 121
rect 55 87 929 93
rect 55 65 929 80
rect 30 40 954 55
<< metal2 >>
rect 18 577 45 580
rect 18 408 21 577
rect 18 3 21 201
rect 30 40 45 540
rect 55 65 70 515
rect 98 478 101 521
rect 170 478 173 580
rect 298 481 301 580
rect 298 478 309 481
rect 138 468 149 471
rect 138 455 141 468
rect 130 448 141 451
rect 130 441 133 448
rect 90 378 93 401
rect 106 258 109 411
rect 138 337 141 448
rect 162 408 165 441
rect 186 408 189 460
rect 218 448 229 451
rect 114 262 118 272
rect 90 168 93 201
rect 114 58 117 262
rect 138 257 141 321
rect 154 315 157 331
rect 186 314 189 331
rect 146 268 149 301
rect 162 132 165 251
rect 18 0 45 3
rect 170 0 173 291
rect 194 138 197 391
rect 218 328 221 448
rect 226 338 229 441
rect 234 418 237 444
rect 250 411 253 461
rect 282 451 285 461
rect 306 448 309 461
rect 234 408 253 411
rect 234 338 237 408
rect 258 348 261 401
rect 202 288 205 321
rect 218 308 221 322
rect 266 311 269 442
rect 298 378 301 441
rect 274 318 277 333
rect 258 308 269 311
rect 218 278 221 301
rect 258 178 261 308
rect 282 268 285 341
rect 290 325 293 361
rect 314 318 317 361
rect 298 298 301 311
rect 322 308 325 464
rect 330 301 333 431
rect 338 398 341 445
rect 354 428 357 465
rect 354 348 357 371
rect 322 298 333 301
rect 282 228 285 247
rect 322 235 325 298
rect 338 247 341 311
rect 346 298 349 321
rect 354 255 357 321
rect 362 278 365 521
rect 426 491 429 580
rect 426 488 453 491
rect 370 408 373 454
rect 394 448 405 451
rect 370 338 373 381
rect 386 378 389 401
rect 378 247 381 301
rect 394 235 397 448
rect 402 398 405 431
rect 410 321 413 471
rect 434 458 437 481
rect 450 461 453 488
rect 466 461 469 471
rect 450 458 461 461
rect 450 451 453 458
rect 434 431 437 441
rect 434 428 445 431
rect 418 348 421 371
rect 426 338 429 381
rect 434 335 437 428
rect 458 381 461 458
rect 458 378 469 381
rect 442 338 445 351
rect 410 318 421 321
rect 418 241 421 318
rect 458 267 461 281
rect 466 261 469 378
rect 474 268 477 330
rect 490 315 493 471
rect 554 461 557 580
rect 530 458 557 461
rect 514 398 517 431
rect 466 258 477 261
rect 498 258 501 351
rect 522 348 525 441
rect 530 388 533 458
rect 538 401 541 454
rect 562 441 565 454
rect 570 451 573 471
rect 578 448 613 451
rect 578 441 581 448
rect 562 438 581 441
rect 554 418 565 421
rect 538 398 549 401
rect 506 338 517 341
rect 506 248 509 338
rect 514 322 517 338
rect 530 328 533 371
rect 538 298 541 334
rect 442 238 445 248
rect 490 245 509 248
rect 362 178 365 231
rect 450 148 453 201
rect 466 138 469 221
rect 482 198 485 241
rect 514 228 517 251
rect 530 218 533 253
rect 546 211 549 398
rect 562 333 565 371
rect 570 338 573 411
rect 578 401 581 431
rect 594 408 597 431
rect 578 398 589 401
rect 610 398 613 448
rect 586 328 589 398
rect 618 351 621 454
rect 666 451 669 461
rect 682 458 685 580
rect 810 478 813 580
rect 882 577 941 580
rect 882 478 885 577
rect 674 441 677 454
rect 690 448 693 461
rect 666 438 677 441
rect 594 319 597 351
rect 610 348 621 351
rect 602 309 605 331
rect 554 268 557 301
rect 554 228 557 244
rect 578 238 581 251
rect 538 208 549 211
rect 298 0 301 101
rect 410 98 413 121
rect 426 0 429 111
rect 538 109 541 208
rect 570 201 573 231
rect 562 198 573 201
rect 562 138 565 198
rect 578 138 581 151
rect 570 118 573 135
rect 586 128 589 264
rect 594 178 597 261
rect 610 178 613 348
rect 618 298 621 321
rect 626 271 629 331
rect 634 325 637 421
rect 658 348 661 361
rect 666 298 669 438
rect 698 378 701 431
rect 714 338 717 451
rect 730 448 733 461
rect 746 428 749 442
rect 770 418 773 451
rect 674 278 677 331
rect 714 301 717 331
rect 722 328 725 371
rect 802 338 805 441
rect 826 378 829 445
rect 826 334 829 351
rect 890 337 893 465
rect 714 298 725 301
rect 722 278 725 298
rect 626 268 637 271
rect 634 257 637 268
rect 658 251 661 261
rect 618 241 622 245
rect 618 238 629 241
rect 602 138 605 151
rect 610 132 614 142
rect 626 138 629 238
rect 634 228 637 241
rect 674 218 677 231
rect 690 211 693 244
rect 698 238 701 257
rect 722 235 725 251
rect 738 247 741 261
rect 690 208 701 211
rect 698 181 701 208
rect 698 178 709 181
rect 554 0 557 111
rect 658 98 661 131
rect 666 118 669 131
rect 682 125 685 151
rect 746 148 749 281
rect 698 121 701 131
rect 682 118 701 121
rect 682 0 685 118
rect 810 0 813 151
rect 882 58 885 301
rect 898 3 901 131
rect 914 65 929 515
rect 939 40 954 540
rect 898 0 941 3
<< metal3 >>
rect 0 517 102 522
rect 361 517 984 522
rect 169 477 222 482
rect 433 477 654 482
rect 737 477 814 482
rect 145 467 470 472
rect 489 467 574 472
rect 177 457 214 462
rect 281 457 310 462
rect 345 457 686 462
rect 137 447 734 452
rect 169 437 230 442
rect 297 437 382 442
rect 401 437 438 442
rect 473 437 566 442
rect 601 437 638 442
rect 721 437 878 442
rect 116 427 278 432
rect 329 427 894 432
rect 233 417 638 422
rect 713 417 774 422
rect 17 407 166 412
rect 185 407 246 412
rect 265 407 494 412
rect 545 407 598 412
rect 0 397 94 402
rect 225 397 342 402
rect 401 397 502 402
rect 513 397 542 402
rect 609 397 984 402
rect 193 387 806 392
rect 217 377 374 382
rect 385 377 430 382
rect 585 377 702 382
rect 737 377 830 382
rect 353 367 726 372
rect 257 357 294 362
rect 313 357 382 362
rect 449 357 662 362
rect 377 352 382 357
rect 97 347 334 352
rect 377 347 502 352
rect 521 347 582 352
rect 593 347 614 352
rect 646 347 830 352
rect 233 337 718 342
rect 153 327 222 332
rect 305 327 462 332
rect 585 327 630 332
rect 641 327 678 332
rect 305 322 310 327
rect 81 317 246 322
rect 273 317 310 322
rect 353 317 774 322
rect 217 307 262 312
rect 273 303 278 317
rect 297 307 878 312
rect 265 302 278 303
rect 217 297 278 302
rect 321 297 350 302
rect 377 297 526 302
rect 537 297 670 302
rect 0 287 984 292
rect 313 277 366 282
rect 457 277 750 282
rect 113 267 150 272
rect 281 267 358 272
rect 473 267 558 272
rect 385 257 470 262
rect 497 257 558 262
rect 593 257 742 262
rect 161 247 374 252
rect 425 247 526 252
rect 561 247 726 252
rect 193 237 254 242
rect 417 237 446 242
rect 537 237 582 242
rect 625 237 702 242
rect 281 227 417 232
rect 513 227 638 232
rect 465 217 678 222
rect 17 197 134 202
rect 481 197 566 202
rect 361 177 446 182
rect 0 167 94 172
rect 979 167 984 172
rect 494 147 606 152
rect 617 147 646 152
rect 681 147 814 152
rect 425 137 510 142
rect 529 137 582 142
rect 609 137 694 142
rect 457 127 702 132
rect 569 117 742 122
rect 401 107 486 112
rect 537 107 558 112
rect 297 97 662 102
rect 0 57 118 62
rect 881 57 984 62
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1490995571
transform 1 0 37 0 1 532
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1490995571
transform 1 0 946 0 1 532
box -7 -7 7 7
use $$M3_M2  $$M3_M2_0
timestamp 1490995571
transform 1 0 100 0 1 520
box -3 -3 3 3
use $$M3_M2  $$M3_M2_1
timestamp 1490995571
transform 1 0 364 0 1 520
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1490995571
transform 1 0 62 0 1 507
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1490995571
transform 1 0 921 0 1 507
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1490995571
transform 1 0 62 0 1 490
box -7 -2 7 2
use $$M3_M2  $$M3_M2_5
timestamp 1490995571
transform 1 0 20 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1490995571
transform 1 0 100 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_7
timestamp 1490995571
transform 1 0 92 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_1
timestamp 1490995571
transform 1 0 148 0 1 470
box -2 -2 2 2
use $$M3_M2  $$M3_M2_2
timestamp 1490995571
transform 1 0 148 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1490995571
transform 1 0 140 0 1 457
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1490995571
transform 1 0 140 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_3
timestamp 1490995571
transform 1 0 132 0 1 443
box -2 -2 2 2
use $$M2_M1  $$M2_M1_4
timestamp 1490995571
transform 1 0 119 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1490995571
transform 1 0 119 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_6
timestamp 1490995571
transform 1 0 108 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_8
timestamp 1490995571
transform 1 0 172 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_5
timestamp 1490995571
transform 1 0 180 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1490995571
transform 1 0 180 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_8
timestamp 1490995571
transform 1 0 188 0 1 459
box -2 -2 2 2
use $$M2_M1  $$M2_M1_9
timestamp 1490995571
transform 1 0 164 0 1 440
box -2 -2 2 2
use $$M2_M1  $$M2_M1_10
timestamp 1490995571
transform 1 0 172 0 1 441
box -2 -2 2 2
use $$M3_M2  $$M3_M2_12
timestamp 1490995571
transform 1 0 172 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_13
timestamp 1490995571
transform 1 0 164 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_16
timestamp 1490995571
transform 1 0 188 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_6
timestamp 1490995571
transform 1 0 220 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_10
timestamp 1490995571
transform 1 0 220 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_7
timestamp 1490995571
transform 1 0 212 0 1 463
box -2 -2 2 2
use $$M3_M2  $$M3_M2_11
timestamp 1490995571
transform 1 0 212 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1490995571
transform 1 0 228 0 1 451
box -2 -2 2 2
use $$M3_M2  $$M3_M2_14
timestamp 1490995571
transform 1 0 228 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_12
timestamp 1490995571
transform 1 0 236 0 1 443
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1490995571
transform 1 0 236 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_18
timestamp 1490995571
transform 1 0 228 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_13
timestamp 1490995571
transform 1 0 252 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_17
timestamp 1490995571
transform 1 0 244 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_19
timestamp 1490995571
transform 1 0 284 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_14
timestamp 1490995571
transform 1 0 284 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_15
timestamp 1490995571
transform 1 0 268 0 1 441
box -2 -2 2 2
use $$M2_M1  $$M2_M1_16
timestamp 1490995571
transform 1 0 276 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_20
timestamp 1490995571
transform 1 0 276 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1490995571
transform 1 0 268 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_17
timestamp 1490995571
transform 1 0 260 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_18
timestamp 1490995571
transform 1 0 308 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_22
timestamp 1490995571
transform 1 0 308 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_22
timestamp 1490995571
transform 1 0 308 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_24
timestamp 1490995571
transform 1 0 300 0 1 441
box -2 -2 2 2
use $$M3_M2  $$M3_M2_24
timestamp 1490995571
transform 1 0 300 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_20
timestamp 1490995571
transform 1 0 324 0 1 463
box -2 -2 2 2
use $$M2_M1  $$M2_M1_21
timestamp 1490995571
transform 1 0 348 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_23
timestamp 1490995571
transform 1 0 348 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_19
timestamp 1490995571
transform 1 0 356 0 1 464
box -2 -2 2 2
use $$M2_M1  $$M2_M1_23
timestamp 1490995571
transform 1 0 340 0 1 443
box -2 -2 2 2
use $$M3_M2  $$M3_M2_25
timestamp 1490995571
transform 1 0 332 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_27
timestamp 1490995571
transform 1 0 340 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_26
timestamp 1490995571
transform 1 0 356 0 1 430
box -3 -3 3 3
use $$M2_M1  $$M2_M1_25
timestamp 1490995571
transform 1 0 372 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_26
timestamp 1490995571
transform 1 0 380 0 1 443
box -2 -2 2 2
use $$M3_M2  $$M3_M2_28
timestamp 1490995571
transform 1 0 380 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_29
timestamp 1490995571
transform 1 0 372 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_27
timestamp 1490995571
transform 1 0 385 0 1 400
box -2 -2 2 2
use $$M3_M2  $$M3_M2_31
timestamp 1490995571
transform 1 0 412 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_29
timestamp 1490995571
transform 1 0 404 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_31
timestamp 1490995571
transform 1 0 404 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_32
timestamp 1490995571
transform 1 0 404 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_32
timestamp 1490995571
transform 1 0 404 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_34
timestamp 1490995571
transform 1 0 404 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_30
timestamp 1490995571
transform 1 0 436 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_28
timestamp 1490995571
transform 1 0 436 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_33
timestamp 1490995571
transform 1 0 436 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_30
timestamp 1490995571
transform 1 0 452 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_33
timestamp 1490995571
transform 1 0 444 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_35
timestamp 1490995571
transform 1 0 468 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_34
timestamp 1490995571
transform 1 0 468 0 1 463
box -2 -2 2 2
use $$M2_M1  $$M2_M1_36
timestamp 1490995571
transform 1 0 476 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_37
timestamp 1490995571
transform 1 0 476 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_36
timestamp 1490995571
transform 1 0 492 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_35
timestamp 1490995571
transform 1 0 492 0 1 450
box -2 -2 2 2
use $$M3_M2  $$M3_M2_39
timestamp 1490995571
transform 1 0 492 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1490995571
transform 1 0 516 0 1 444
box -2 -2 2 2
use $$M3_M2  $$M3_M2_38
timestamp 1490995571
transform 1 0 516 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_38
timestamp 1490995571
transform 1 0 524 0 1 440
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1490995571
transform 1 0 516 0 1 430
box -2 -2 2 2
use $$M2_M1  $$M2_M1_40
timestamp 1490995571
transform 1 0 500 0 1 400
box -2 -2 2 2
use $$M3_M2  $$M3_M2_40
timestamp 1490995571
transform 1 0 500 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_41
timestamp 1490995571
transform 1 0 516 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_41
timestamp 1490995571
transform 1 0 540 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1490995571
transform 1 0 572 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1490995571
transform 1 0 564 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_45
timestamp 1490995571
transform 1 0 572 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_45
timestamp 1490995571
transform 1 0 564 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_42
timestamp 1490995571
transform 1 0 556 0 1 420
box -2 -2 2 2
use $$M3_M2  $$M3_M2_46
timestamp 1490995571
transform 1 0 564 0 1 420
box -3 -3 3 3
use $$M2_M1  $$M2_M1_43
timestamp 1490995571
transform 1 0 548 0 1 410
box -2 -2 2 2
use $$M3_M2  $$M3_M2_42
timestamp 1490995571
transform 1 0 548 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_43
timestamp 1490995571
transform 1 0 540 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_47
timestamp 1490995571
transform 1 0 572 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_46
timestamp 1490995571
transform 1 0 580 0 1 430
box -2 -2 2 2
use $$M2_M1  $$M2_M1_47
timestamp 1490995571
transform 1 0 612 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_48
timestamp 1490995571
transform 1 0 620 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1490995571
transform 1 0 604 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1490995571
transform 1 0 604 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_50
timestamp 1490995571
transform 1 0 596 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_49
timestamp 1490995571
transform 1 0 596 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_50
timestamp 1490995571
transform 1 0 612 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_51
timestamp 1490995571
transform 1 0 652 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_51
timestamp 1490995571
transform 1 0 652 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_52
timestamp 1490995571
transform 1 0 636 0 1 443
box -2 -2 2 2
use $$M3_M2  $$M3_M2_52
timestamp 1490995571
transform 1 0 636 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_53
timestamp 1490995571
transform 1 0 636 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_54
timestamp 1490995571
transform 1 0 668 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1490995571
transform 1 0 668 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_55
timestamp 1490995571
transform 1 0 676 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_55
timestamp 1490995571
transform 1 0 684 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_53
timestamp 1490995571
transform 1 0 692 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_56
timestamp 1490995571
transform 1 0 692 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_63
timestamp 1490995571
transform 1 0 700 0 1 430
box -2 -2 2 2
use $$M2_M1  $$M2_M1_56
timestamp 1490995571
transform 1 0 716 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_57
timestamp 1490995571
transform 1 0 740 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_57
timestamp 1490995571
transform 1 0 740 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_58
timestamp 1490995571
transform 1 0 732 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1490995571
transform 1 0 732 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_62
timestamp 1490995571
transform 1 0 724 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_60
timestamp 1490995571
transform 1 0 724 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_61
timestamp 1490995571
transform 1 0 716 0 1 420
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1490995571
transform 1 0 748 0 1 441
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1490995571
transform 1 0 748 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_58
timestamp 1490995571
transform 1 0 812 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1490995571
transform 1 0 772 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_60
timestamp 1490995571
transform 1 0 828 0 1 444
box -2 -2 2 2
use $$M2_M1  $$M2_M1_64
timestamp 1490995571
transform 1 0 804 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1490995571
transform 1 0 772 0 1 420
box -3 -3 3 3
use $$M2_M1  $$M2_M1_65
timestamp 1490995571
transform 1 0 884 0 1 480
box -2 -2 2 2
use $$M2_M1  $$M2_M1_67
timestamp 1490995571
transform 1 0 876 0 1 441
box -2 -2 2 2
use $$M3_M2  $$M3_M2_64
timestamp 1490995571
transform 1 0 876 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_66
timestamp 1490995571
transform 1 0 892 0 1 464
box -2 -2 2 2
use $$M3_M2  $$M3_M2_65
timestamp 1490995571
transform 1 0 892 0 1 430
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1490995571
transform 1 0 921 0 1 490
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1490995571
transform 1 0 37 0 1 390
box -7 -2 7 2
use FILL  FILL_0
timestamp 1490995571
transform 1 0 80 0 -1 490
box -8 -3 16 105
use FILL  FILL_1
timestamp 1490995571
transform 1 0 88 0 -1 490
box -8 -3 16 105
use FILL  FILL_2
timestamp 1490995571
transform 1 0 96 0 -1 490
box -8 -3 16 105
use FILL  FILL_3
timestamp 1490995571
transform 1 0 104 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1490995571
transform -1 0 144 0 -1 490
box -8 -3 34 105
use FILL  FILL_4
timestamp 1490995571
transform 1 0 144 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1490995571
transform 1 0 152 0 -1 490
box -8 -3 32 105
use $$M3_M2  $$M3_M2_66
timestamp 1490995571
transform 1 0 196 0 1 390
box -3 -3 3 3
use INVX2  INVX2_0
timestamp 1490995571
transform -1 0 192 0 -1 490
box -9 -3 26 105
use FILL  FILL_5
timestamp 1490995571
transform 1 0 192 0 -1 490
box -8 -3 16 105
use FILL  FILL_6
timestamp 1490995571
transform 1 0 200 0 -1 490
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1490995571
transform -1 0 240 0 -1 490
box -7 -3 39 105
use FILL  FILL_7
timestamp 1490995571
transform 1 0 240 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1490995571
transform 1 0 248 0 -1 490
box -8 -3 32 105
use INVX2  INVX2_1
timestamp 1490995571
transform -1 0 288 0 -1 490
box -9 -3 26 105
use FILL  FILL_8
timestamp 1490995571
transform 1 0 288 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1490995571
transform -1 0 320 0 -1 490
box -8 -3 32 105
use FILL  FILL_9
timestamp 1490995571
transform 1 0 320 0 -1 490
box -8 -3 16 105
use FILL  FILL_10
timestamp 1490995571
transform 1 0 328 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1490995571
transform -1 0 360 0 -1 490
box -8 -3 32 105
use FILL  FILL_11
timestamp 1490995571
transform 1 0 360 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1490995571
transform 1 0 368 0 -1 490
box -8 -3 34 105
use FILL  FILL_12
timestamp 1490995571
transform 1 0 400 0 -1 490
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1490995571
transform -1 0 432 0 -1 490
box -8 -3 32 105
use FILL  FILL_13
timestamp 1490995571
transform 1 0 432 0 -1 490
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1490995571
transform -1 0 456 0 -1 490
box -9 -3 26 105
use FILL  FILL_14
timestamp 1490995571
transform 1 0 456 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1490995571
transform 1 0 464 0 -1 490
box -8 -3 32 105
use FILL  FILL_15
timestamp 1490995571
transform 1 0 488 0 -1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_67
timestamp 1490995571
transform 1 0 532 0 1 390
box -3 -3 3 3
use NAND3X1  NAND3X1_0
timestamp 1490995571
transform -1 0 528 0 -1 490
box -8 -3 40 105
use FILL  FILL_16
timestamp 1490995571
transform 1 0 528 0 -1 490
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1490995571
transform 1 0 536 0 -1 490
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1490995571
transform -1 0 568 0 -1 490
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1490995571
transform 1 0 568 0 -1 490
box -9 -3 26 105
use FILL  FILL_17
timestamp 1490995571
transform 1 0 584 0 -1 490
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1490995571
transform -1 0 616 0 -1 490
box -8 -3 32 105
use FILL  FILL_18
timestamp 1490995571
transform 1 0 616 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1490995571
transform 1 0 624 0 -1 490
box -8 -3 34 105
use INVX2  INVX2_6
timestamp 1490995571
transform -1 0 672 0 -1 490
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1490995571
transform 1 0 672 0 -1 490
box -9 -3 26 105
use FILL  FILL_19
timestamp 1490995571
transform 1 0 688 0 -1 490
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1490995571
transform -1 0 720 0 -1 490
box -8 -3 32 105
use FILL  FILL_20
timestamp 1490995571
transform 1 0 720 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1490995571
transform 1 0 728 0 -1 490
box -8 -3 32 105
use FILL  FILL_21
timestamp 1490995571
transform 1 0 752 0 -1 490
box -8 -3 16 105
use FILL  FILL_22
timestamp 1490995571
transform 1 0 760 0 -1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_68
timestamp 1490995571
transform 1 0 804 0 1 390
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_0
timestamp 1490995571
transform -1 0 864 0 -1 490
box -8 -3 104 105
use FILL  FILL_23
timestamp 1490995571
transform 1 0 864 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1490995571
transform -1 0 896 0 -1 490
box -8 -3 32 105
use FILL  FILL_24
timestamp 1490995571
transform 1 0 896 0 -1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1490995571
transform 1 0 946 0 1 390
box -7 -2 7 2
use $$M2_M1  $$M2_M1_68
timestamp 1490995571
transform 1 0 92 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_69
timestamp 1490995571
transform 1 0 100 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_69
timestamp 1490995571
transform 1 0 100 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_70
timestamp 1490995571
transform 1 0 84 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_70
timestamp 1490995571
transform 1 0 84 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_71
timestamp 1490995571
transform 1 0 140 0 1 339
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1490995571
transform 1 0 140 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_71
timestamp 1490995571
transform 1 0 156 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_72
timestamp 1490995571
transform 1 0 156 0 1 317
box -2 -2 2 2
use $$M2_M1  $$M2_M1_73
timestamp 1490995571
transform 1 0 148 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_73
timestamp 1490995571
transform 1 0 188 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_75
timestamp 1490995571
transform 1 0 188 0 1 316
box -2 -2 2 2
use $$M2_M1  $$M2_M1_74
timestamp 1490995571
transform 1 0 204 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_74
timestamp 1490995571
transform 1 0 220 0 1 380
box -3 -3 3 3
use $$M2_M1  $$M2_M1_76
timestamp 1490995571
transform 1 0 236 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_77
timestamp 1490995571
transform 1 0 228 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_76
timestamp 1490995571
transform 1 0 220 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_78
timestamp 1490995571
transform 1 0 220 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_82
timestamp 1490995571
transform 1 0 220 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_83
timestamp 1490995571
transform 1 0 220 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_75
timestamp 1490995571
transform 1 0 236 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_82
timestamp 1490995571
transform 1 0 244 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_80
timestamp 1490995571
transform 1 0 244 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_77
timestamp 1490995571
transform 1 0 260 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_79
timestamp 1490995571
transform 1 0 260 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_79
timestamp 1490995571
transform 1 0 292 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_80
timestamp 1490995571
transform 1 0 284 0 1 340
box -2 -2 2 2
use $$M2_M1  $$M2_M1_81
timestamp 1490995571
transform 1 0 276 0 1 331
box -2 -2 2 2
use $$M3_M2  $$M3_M2_81
timestamp 1490995571
transform 1 0 276 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_84
timestamp 1490995571
transform 1 0 260 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_83
timestamp 1490995571
transform 1 0 292 0 1 327
box -2 -2 2 2
use $$M3_M2  $$M3_M2_78
timestamp 1490995571
transform 1 0 300 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_85
timestamp 1490995571
transform 1 0 316 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_84
timestamp 1490995571
transform 1 0 308 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_86
timestamp 1490995571
transform 1 0 308 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_87
timestamp 1490995571
transform 1 0 300 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_86
timestamp 1490995571
transform 1 0 300 0 1 300
box -2 -2 2 2
use $$M2_M1  $$M2_M1_85
timestamp 1490995571
transform 1 0 316 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_93
timestamp 1490995571
transform 1 0 332 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_88
timestamp 1490995571
transform 1 0 324 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_89
timestamp 1490995571
transform 1 0 324 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_90
timestamp 1490995571
transform 1 0 372 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_92
timestamp 1490995571
transform 1 0 356 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_87
timestamp 1490995571
transform 1 0 356 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_91
timestamp 1490995571
transform 1 0 388 0 1 380
box -3 -3 3 3
use $$M2_M1  $$M2_M1_88
timestamp 1490995571
transform 1 0 380 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_94
timestamp 1490995571
transform 1 0 380 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_89
timestamp 1490995571
transform 1 0 372 0 1 340
box -2 -2 2 2
use $$M2_M1  $$M2_M1_91
timestamp 1490995571
transform 1 0 348 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_96
timestamp 1490995571
transform 1 0 340 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_90
timestamp 1490995571
transform 1 0 356 0 1 323
box -2 -2 2 2
use $$M3_M2  $$M3_M2_95
timestamp 1490995571
transform 1 0 356 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_97
timestamp 1490995571
transform 1 0 348 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_92
timestamp 1490995571
transform 1 0 388 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_98
timestamp 1490995571
transform 1 0 388 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_99
timestamp 1490995571
transform 1 0 380 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_100
timestamp 1490995571
transform 1 0 428 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_101
timestamp 1490995571
transform 1 0 420 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_94
timestamp 1490995571
transform 1 0 420 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_96
timestamp 1490995571
transform 1 0 412 0 1 320
box -2 -2 2 2
use $$M2_M1  $$M2_M1_93
timestamp 1490995571
transform 1 0 452 0 1 360
box -2 -2 2 2
use $$M3_M2  $$M3_M2_102
timestamp 1490995571
transform 1 0 452 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_95
timestamp 1490995571
transform 1 0 444 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_97
timestamp 1490995571
transform 1 0 428 0 1 340
box -2 -2 2 2
use $$M2_M1  $$M2_M1_98
timestamp 1490995571
transform 1 0 436 0 1 337
box -2 -2 2 2
use $$M3_M2  $$M3_M2_103
timestamp 1490995571
transform 1 0 444 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_99
timestamp 1490995571
transform 1 0 460 0 1 333
box -2 -2 2 2
use $$M3_M2  $$M3_M2_104
timestamp 1490995571
transform 1 0 460 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_100
timestamp 1490995571
transform 1 0 476 0 1 329
box -2 -2 2 2
use $$M3_M2  $$M3_M2_106
timestamp 1490995571
transform 1 0 500 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_101
timestamp 1490995571
transform 1 0 492 0 1 317
box -2 -2 2 2
use $$M3_M2  $$M3_M2_105
timestamp 1490995571
transform 1 0 532 0 1 370
box -3 -3 3 3
use $$M3_M2  $$M3_M2_107
timestamp 1490995571
transform 1 0 524 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_108
timestamp 1490995571
transform 1 0 516 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_109
timestamp 1490995571
transform 1 0 564 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_102
timestamp 1490995571
transform 1 0 556 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_111
timestamp 1490995571
transform 1 0 556 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_110
timestamp 1490995571
transform 1 0 588 0 1 380
box -3 -3 3 3
use $$M2_M1  $$M2_M1_103
timestamp 1490995571
transform 1 0 580 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_112
timestamp 1490995571
transform 1 0 580 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_104
timestamp 1490995571
transform 1 0 572 0 1 340
box -2 -2 2 2
use $$M2_M1  $$M2_M1_107
timestamp 1490995571
transform 1 0 532 0 1 330
box -2 -2 2 2
use $$M2_M1  $$M2_M1_106
timestamp 1490995571
transform 1 0 540 0 1 333
box -2 -2 2 2
use $$M2_M1  $$M2_M1_105
timestamp 1490995571
transform 1 0 564 0 1 335
box -2 -2 2 2
use $$M2_M1  $$M2_M1_108
timestamp 1490995571
transform 1 0 516 0 1 324
box -2 -2 2 2
use $$M2_M1  $$M2_M1_109
timestamp 1490995571
transform 1 0 524 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_113
timestamp 1490995571
transform 1 0 524 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_114
timestamp 1490995571
transform 1 0 540 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_110
timestamp 1490995571
transform 1 0 556 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_115
timestamp 1490995571
transform 1 0 596 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_116
timestamp 1490995571
transform 1 0 612 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_118
timestamp 1490995571
transform 1 0 588 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_119
timestamp 1490995571
transform 1 0 604 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_112
timestamp 1490995571
transform 1 0 596 0 1 321
box -2 -2 2 2
use $$M2_M1  $$M2_M1_118
timestamp 1490995571
transform 1 0 604 0 1 311
box -2 -2 2 2
use $$M2_M1  $$M2_M1_111
timestamp 1490995571
transform 1 0 620 0 1 339
box -2 -2 2 2
use $$M3_M2  $$M3_M2_117
timestamp 1490995571
transform 1 0 620 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_122
timestamp 1490995571
transform 1 0 628 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_120
timestamp 1490995571
transform 1 0 660 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_113
timestamp 1490995571
transform 1 0 649 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_121
timestamp 1490995571
transform 1 0 649 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_114
timestamp 1490995571
transform 1 0 660 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_117
timestamp 1490995571
transform 1 0 620 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_127
timestamp 1490995571
transform 1 0 620 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_119
timestamp 1490995571
transform 1 0 636 0 1 327
box -2 -2 2 2
use $$M2_M1  $$M2_M1_115
timestamp 1490995571
transform 1 0 644 0 1 331
box -2 -2 2 2
use $$M3_M2  $$M3_M2_123
timestamp 1490995571
transform 1 0 644 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_126
timestamp 1490995571
transform 1 0 676 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_129
timestamp 1490995571
transform 1 0 668 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_124
timestamp 1490995571
transform 1 0 700 0 1 380
box -3 -3 3 3
use $$M2_M1  $$M2_M1_116
timestamp 1490995571
transform 1 0 700 0 1 370
box -2 -2 2 2
use $$M3_M2  $$M3_M2_125
timestamp 1490995571
transform 1 0 700 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_120
timestamp 1490995571
transform 1 0 692 0 1 322
box -2 -2 2 2
use $$M3_M2  $$M3_M2_128
timestamp 1490995571
transform 1 0 692 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_121
timestamp 1490995571
transform 1 0 740 0 1 380
box -2 -2 2 2
use $$M3_M2  $$M3_M2_130
timestamp 1490995571
transform 1 0 740 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_131
timestamp 1490995571
transform 1 0 724 0 1 370
box -3 -3 3 3
use $$M3_M2  $$M3_M2_132
timestamp 1490995571
transform 1 0 716 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_122
timestamp 1490995571
transform 1 0 716 0 1 330
box -2 -2 2 2
use $$M2_M1  $$M2_M1_123
timestamp 1490995571
transform 1 0 724 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_133
timestamp 1490995571
transform 1 0 828 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_134
timestamp 1490995571
transform 1 0 828 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_124
timestamp 1490995571
transform 1 0 804 0 1 340
box -2 -2 2 2
use $$M2_M1  $$M2_M1_125
timestamp 1490995571
transform 1 0 828 0 1 336
box -2 -2 2 2
use $$M2_M1  $$M2_M1_126
timestamp 1490995571
transform 1 0 772 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_135
timestamp 1490995571
transform 1 0 772 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_170
timestamp 1490995571
transform 1 0 876 0 1 311
box -2 -2 2 2
use $$M3_M2  $$M3_M2_177
timestamp 1490995571
transform 1 0 876 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_169
timestamp 1490995571
transform 1 0 892 0 1 339
box -2 -2 2 2
use $$M2_M1  $$M2_M1_171
timestamp 1490995571
transform 1 0 884 0 1 300
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1490995571
transform 1 0 62 0 1 290
box -7 -2 7 2
use NAND2X1  NAND2X1_3
timestamp 1490995571
transform 1 0 80 0 1 290
box -8 -3 32 105
use FILL  FILL_25
timestamp 1490995571
transform -1 0 112 0 1 290
box -8 -3 16 105
use FILL  FILL_27
timestamp 1490995571
transform -1 0 120 0 1 290
box -8 -3 16 105
use FILL  FILL_28
timestamp 1490995571
transform -1 0 128 0 1 290
box -8 -3 16 105
use FILL  FILL_29
timestamp 1490995571
transform -1 0 136 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1490995571
transform -1 0 160 0 1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_136
timestamp 1490995571
transform 1 0 172 0 1 290
box -3 -3 3 3
use FILL  FILL_30
timestamp 1490995571
transform -1 0 168 0 1 290
box -8 -3 16 105
use FILL  FILL_31
timestamp 1490995571
transform -1 0 176 0 1 290
box -8 -3 16 105
use FILL  FILL_32
timestamp 1490995571
transform -1 0 184 0 1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_137
timestamp 1490995571
transform 1 0 204 0 1 290
box -3 -3 3 3
use NOR2X1  NOR2X1_8
timestamp 1490995571
transform 1 0 184 0 1 290
box -8 -3 32 105
use FILL  FILL_33
timestamp 1490995571
transform -1 0 216 0 1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1490995571
transform 1 0 216 0 1 290
box -8 -3 32 105
use FILL  FILL_44
timestamp 1490995571
transform -1 0 248 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1490995571
transform -1 0 280 0 1 290
box -8 -3 40 105
use FILL  FILL_45
timestamp 1490995571
transform -1 0 288 0 1 290
box -8 -3 16 105
use INVX2  INVX2_8
timestamp 1490995571
transform 1 0 288 0 1 290
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1490995571
transform 1 0 304 0 1 290
box -9 -3 26 105
use FILL  FILL_47
timestamp 1490995571
transform -1 0 328 0 1 290
box -8 -3 16 105
use FILL  FILL_48
timestamp 1490995571
transform -1 0 336 0 1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1490995571
transform 1 0 336 0 1 290
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1490995571
transform 1 0 360 0 1 290
box -8 -3 32 105
use FILL  FILL_50
timestamp 1490995571
transform -1 0 392 0 1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1490995571
transform 1 0 392 0 1 290
box -8 -3 32 105
use FILL  FILL_52
timestamp 1490995571
transform -1 0 424 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1490995571
transform 1 0 424 0 1 290
box -8 -3 40 105
use FILL  FILL_54
timestamp 1490995571
transform -1 0 464 0 1 290
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1490995571
transform 1 0 464 0 1 290
box -7 -3 39 105
use FILL  FILL_57
timestamp 1490995571
transform -1 0 504 0 1 290
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1490995571
transform 1 0 504 0 1 290
box -8 -3 46 105
use NAND3X1  NAND3X1_3
timestamp 1490995571
transform -1 0 576 0 1 290
box -8 -3 40 105
use FILL  FILL_58
timestamp 1490995571
transform -1 0 584 0 1 290
box -8 -3 16 105
use INVX2  INVX2_10
timestamp 1490995571
transform -1 0 600 0 1 290
box -9 -3 26 105
use NOR2X1  NOR2X1_9
timestamp 1490995571
transform 1 0 600 0 1 290
box -8 -3 32 105
use FILL  FILL_61
timestamp 1490995571
transform -1 0 632 0 1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1490995571
transform 1 0 632 0 1 290
box -8 -3 34 105
use FILL  FILL_64
timestamp 1490995571
transform -1 0 672 0 1 290
box -8 -3 16 105
use FILL  FILL_65
timestamp 1490995571
transform -1 0 680 0 1 290
box -8 -3 16 105
use FILL  FILL_66
timestamp 1490995571
transform -1 0 688 0 1 290
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1490995571
transform 1 0 688 0 1 290
box -9 -3 26 105
use FILL  FILL_67
timestamp 1490995571
transform -1 0 712 0 1 290
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1490995571
transform 1 0 712 0 1 290
box -8 -3 40 105
use FILL  FILL_70
timestamp 1490995571
transform -1 0 752 0 1 290
box -8 -3 16 105
use FILL  FILL_71
timestamp 1490995571
transform -1 0 760 0 1 290
box -8 -3 16 105
use FILL  FILL_72
timestamp 1490995571
transform -1 0 768 0 1 290
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_2
timestamp 1490995571
transform -1 0 864 0 1 290
box -8 -3 104 105
use FILL  FILL_73
timestamp 1490995571
transform -1 0 872 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1490995571
transform 1 0 872 0 1 290
box -8 -3 32 105
use FILL  FILL_74
timestamp 1490995571
transform -1 0 904 0 1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_6
timestamp 1490995571
transform 1 0 921 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_139
timestamp 1490995571
transform 1 0 20 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_138
timestamp 1490995571
transform 1 0 116 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_127
timestamp 1490995571
transform 1 0 116 0 1 264
box -2 -2 2 2
use $$M2_M1  $$M2_M1_128
timestamp 1490995571
transform 1 0 108 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_129
timestamp 1490995571
transform 1 0 92 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_140
timestamp 1490995571
transform 1 0 148 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_130
timestamp 1490995571
transform 1 0 140 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_135
timestamp 1490995571
transform 1 0 132 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_146
timestamp 1490995571
transform 1 0 132 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_143
timestamp 1490995571
transform 1 0 164 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_144
timestamp 1490995571
transform 1 0 196 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_131
timestamp 1490995571
transform 1 0 220 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_132
timestamp 1490995571
transform 1 0 316 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_141
timestamp 1490995571
transform 1 0 316 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_142
timestamp 1490995571
transform 1 0 284 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_133
timestamp 1490995571
transform 1 0 284 0 1 246
box -2 -2 2 2
use $$M2_M1  $$M2_M1_134
timestamp 1490995571
transform 1 0 252 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_145
timestamp 1490995571
transform 1 0 252 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_147
timestamp 1490995571
transform 1 0 284 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_149
timestamp 1490995571
transform 1 0 364 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_148
timestamp 1490995571
transform 1 0 356 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_136
timestamp 1490995571
transform 1 0 356 0 1 257
box -2 -2 2 2
use $$M2_M1  $$M2_M1_137
timestamp 1490995571
transform 1 0 340 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_138
timestamp 1490995571
transform 1 0 324 0 1 237
box -2 -2 2 2
use $$M3_M2  $$M3_M2_150
timestamp 1490995571
transform 1 0 388 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_139
timestamp 1490995571
transform 1 0 388 0 1 257
box -2 -2 2 2
use $$M2_M1  $$M2_M1_140
timestamp 1490995571
transform 1 0 372 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_151
timestamp 1490995571
transform 1 0 372 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_141
timestamp 1490995571
transform 1 0 380 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_143
timestamp 1490995571
transform 1 0 364 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_142
timestamp 1490995571
transform 1 0 396 0 1 237
box -2 -2 2 2
use $$M2_M1  $$M2_M1_144
timestamp 1490995571
transform 1 0 428 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_152
timestamp 1490995571
transform 1 0 428 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_145
timestamp 1490995571
transform 1 0 420 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_153
timestamp 1490995571
transform 1 0 420 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_146
timestamp 1490995571
transform 1 0 415 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_154
timestamp 1490995571
transform 1 0 415 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_149
timestamp 1490995571
transform 1 0 444 0 1 247
box -2 -2 2 2
use $$M3_M2  $$M3_M2_159
timestamp 1490995571
transform 1 0 444 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_155
timestamp 1490995571
transform 1 0 460 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_147
timestamp 1490995571
transform 1 0 460 0 1 269
box -2 -2 2 2
use $$M2_M1  $$M2_M1_152
timestamp 1490995571
transform 1 0 452 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_156
timestamp 1490995571
transform 1 0 476 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_157
timestamp 1490995571
transform 1 0 468 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_148
timestamp 1490995571
transform 1 0 476 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_160
timestamp 1490995571
transform 1 0 468 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_158
timestamp 1490995571
transform 1 0 500 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_150
timestamp 1490995571
transform 1 0 492 0 1 247
box -2 -2 2 2
use $$M2_M1  $$M2_M1_151
timestamp 1490995571
transform 1 0 484 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_161
timestamp 1490995571
transform 1 0 484 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_154
timestamp 1490995571
transform 1 0 516 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_155
timestamp 1490995571
transform 1 0 524 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_153
timestamp 1490995571
transform 1 0 532 0 1 252
box -2 -2 2 2
use $$M3_M2  $$M3_M2_162
timestamp 1490995571
transform 1 0 524 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_163
timestamp 1490995571
transform 1 0 556 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_164
timestamp 1490995571
transform 1 0 556 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_156
timestamp 1490995571
transform 1 0 556 0 1 257
box -2 -2 2 2
use $$M2_M1  $$M2_M1_157
timestamp 1490995571
transform 1 0 564 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_165
timestamp 1490995571
transform 1 0 564 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_159
timestamp 1490995571
transform 1 0 540 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_166
timestamp 1490995571
transform 1 0 540 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_158
timestamp 1490995571
transform 1 0 556 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_167
timestamp 1490995571
transform 1 0 516 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_168
timestamp 1490995571
transform 1 0 532 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_169
timestamp 1490995571
transform 1 0 556 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_161
timestamp 1490995571
transform 1 0 588 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_171
timestamp 1490995571
transform 1 0 596 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_162
timestamp 1490995571
transform 1 0 580 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_172
timestamp 1490995571
transform 1 0 580 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_160
timestamp 1490995571
transform 1 0 572 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_170
timestamp 1490995571
transform 1 0 564 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_164
timestamp 1490995571
transform 1 0 620 0 1 244
box -2 -2 2 2
use $$M2_M1  $$M2_M1_163
timestamp 1490995571
transform 1 0 636 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_166
timestamp 1490995571
transform 1 0 612 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_173
timestamp 1490995571
transform 1 0 628 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_165
timestamp 1490995571
transform 1 0 636 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_174
timestamp 1490995571
transform 1 0 636 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_175
timestamp 1490995571
transform 1 0 660 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_167
timestamp 1490995571
transform 1 0 660 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_168
timestamp 1490995571
transform 1 0 652 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_176
timestamp 1490995571
transform 1 0 652 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_172
timestamp 1490995571
transform 1 0 676 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_173
timestamp 1490995571
transform 1 0 700 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_174
timestamp 1490995571
transform 1 0 692 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_175
timestamp 1490995571
transform 1 0 676 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_179
timestamp 1490995571
transform 1 0 676 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_178
timestamp 1490995571
transform 1 0 700 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_176
timestamp 1490995571
transform 1 0 724 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_180
timestamp 1490995571
transform 1 0 748 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_181
timestamp 1490995571
transform 1 0 740 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_182
timestamp 1490995571
transform 1 0 724 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_177
timestamp 1490995571
transform 1 0 748 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_178
timestamp 1490995571
transform 1 0 740 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_179
timestamp 1490995571
transform 1 0 724 0 1 237
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1490995571
transform 1 0 37 0 1 190
box -7 -2 7 2
use FILL  FILL_26
timestamp 1490995571
transform 1 0 80 0 -1 290
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1490995571
transform -1 0 120 0 -1 290
box -8 -3 40 105
use FILL  FILL_34
timestamp 1490995571
transform 1 0 120 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1490995571
transform -1 0 144 0 -1 290
box -9 -3 26 105
use FILL  FILL_35
timestamp 1490995571
transform 1 0 144 0 -1 290
box -8 -3 16 105
use FILL  FILL_36
timestamp 1490995571
transform 1 0 152 0 -1 290
box -8 -3 16 105
use FILL  FILL_37
timestamp 1490995571
transform 1 0 160 0 -1 290
box -8 -3 16 105
use FILL  FILL_38
timestamp 1490995571
transform 1 0 168 0 -1 290
box -8 -3 16 105
use FILL  FILL_39
timestamp 1490995571
transform 1 0 176 0 -1 290
box -8 -3 16 105
use FILL  FILL_40
timestamp 1490995571
transform 1 0 184 0 -1 290
box -8 -3 16 105
use FILL  FILL_41
timestamp 1490995571
transform 1 0 192 0 -1 290
box -8 -3 16 105
use FILL  FILL_42
timestamp 1490995571
transform 1 0 200 0 -1 290
box -8 -3 16 105
use FILL  FILL_43
timestamp 1490995571
transform 1 0 208 0 -1 290
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_1
timestamp 1490995571
transform -1 0 312 0 -1 290
box -8 -3 104 105
use FILL  FILL_46
timestamp 1490995571
transform 1 0 312 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1490995571
transform -1 0 352 0 -1 290
box -8 -3 34 105
use FILL  FILL_49
timestamp 1490995571
transform 1 0 352 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1490995571
transform -1 0 392 0 -1 290
box -8 -3 34 105
use FILL  FILL_51
timestamp 1490995571
transform 1 0 392 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1490995571
transform -1 0 432 0 -1 290
box -8 -3 34 105
use FILL  FILL_53
timestamp 1490995571
transform 1 0 432 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1490995571
transform -1 0 464 0 -1 290
box -8 -3 32 105
use FILL  FILL_55
timestamp 1490995571
transform 1 0 464 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1490995571
transform 1 0 472 0 -1 290
box -8 -3 32 105
use FILL  FILL_56
timestamp 1490995571
transform 1 0 496 0 -1 290
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1490995571
transform -1 0 544 0 -1 290
box -8 -3 46 105
use OAI21X1  OAI21X1_7
timestamp 1490995571
transform 1 0 544 0 -1 290
box -8 -3 34 105
use FILL  FILL_59
timestamp 1490995571
transform 1 0 576 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1490995571
transform 1 0 584 0 -1 290
box -8 -3 32 105
use FILL  FILL_60
timestamp 1490995571
transform 1 0 608 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1490995571
transform -1 0 640 0 -1 290
box -8 -3 32 105
use FILL  FILL_62
timestamp 1490995571
transform 1 0 640 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_13
timestamp 1490995571
transform -1 0 664 0 -1 290
box -9 -3 26 105
use FILL  FILL_63
timestamp 1490995571
transform 1 0 664 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1490995571
transform -1 0 704 0 -1 290
box -8 -3 34 105
use FILL  FILL_68
timestamp 1490995571
transform 1 0 704 0 -1 290
box -8 -3 16 105
use FILL  FILL_69
timestamp 1490995571
transform 1 0 712 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1490995571
transform -1 0 752 0 -1 290
box -8 -3 34 105
use FILL  FILL_75
timestamp 1490995571
transform 1 0 752 0 -1 290
box -8 -3 16 105
use FILL  FILL_76
timestamp 1490995571
transform 1 0 760 0 -1 290
box -8 -3 16 105
use FILL  FILL_77
timestamp 1490995571
transform 1 0 768 0 -1 290
box -8 -3 16 105
use FILL  FILL_78
timestamp 1490995571
transform 1 0 776 0 -1 290
box -8 -3 16 105
use FILL  FILL_79
timestamp 1490995571
transform 1 0 784 0 -1 290
box -8 -3 16 105
use FILL  FILL_80
timestamp 1490995571
transform 1 0 792 0 -1 290
box -8 -3 16 105
use FILL  FILL_81
timestamp 1490995571
transform 1 0 800 0 -1 290
box -8 -3 16 105
use FILL  FILL_82
timestamp 1490995571
transform 1 0 808 0 -1 290
box -8 -3 16 105
use FILL  FILL_83
timestamp 1490995571
transform 1 0 816 0 -1 290
box -8 -3 16 105
use FILL  FILL_84
timestamp 1490995571
transform 1 0 824 0 -1 290
box -8 -3 16 105
use FILL  FILL_85
timestamp 1490995571
transform 1 0 832 0 -1 290
box -8 -3 16 105
use FILL  FILL_86
timestamp 1490995571
transform 1 0 840 0 -1 290
box -8 -3 16 105
use FILL  FILL_87
timestamp 1490995571
transform 1 0 848 0 -1 290
box -8 -3 16 105
use FILL  FILL_88
timestamp 1490995571
transform 1 0 856 0 -1 290
box -8 -3 16 105
use FILL  FILL_89
timestamp 1490995571
transform 1 0 864 0 -1 290
box -8 -3 16 105
use FILL  FILL_90
timestamp 1490995571
transform 1 0 872 0 -1 290
box -8 -3 16 105
use FILL  FILL_91
timestamp 1490995571
transform 1 0 880 0 -1 290
box -8 -3 16 105
use FILL  FILL_92
timestamp 1490995571
transform 1 0 888 0 -1 290
box -8 -3 16 105
use FILL  FILL_93
timestamp 1490995571
transform 1 0 896 0 -1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_7
timestamp 1490995571
transform 1 0 946 0 1 190
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_8
timestamp 1490995571
transform 1 0 62 0 1 90
box -7 -2 7 2
use $$M3_M2  $$M3_M2_183
timestamp 1490995571
transform 1 0 92 0 1 170
box -3 -3 3 3
use FILL  FILL_94
timestamp 1490995571
transform -1 0 88 0 1 90
box -8 -3 16 105
use FILL  FILL_95
timestamp 1490995571
transform -1 0 96 0 1 90
box -8 -3 16 105
use FILL  FILL_96
timestamp 1490995571
transform -1 0 104 0 1 90
box -8 -3 16 105
use FILL  FILL_97
timestamp 1490995571
transform -1 0 112 0 1 90
box -8 -3 16 105
use FILL  FILL_98
timestamp 1490995571
transform -1 0 120 0 1 90
box -8 -3 16 105
use FILL  FILL_99
timestamp 1490995571
transform -1 0 128 0 1 90
box -8 -3 16 105
use FILL  FILL_100
timestamp 1490995571
transform -1 0 136 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_181
timestamp 1490995571
transform 1 0 196 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_182
timestamp 1490995571
transform 1 0 164 0 1 134
box -2 -2 2 2
use DFFPOSX1  DFFPOSX1_3
timestamp 1490995571
transform 1 0 136 0 1 90
box -8 -3 104 105
use FILL  FILL_101
timestamp 1490995571
transform -1 0 240 0 1 90
box -8 -3 16 105
use FILL  FILL_102
timestamp 1490995571
transform -1 0 248 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_180
timestamp 1490995571
transform 1 0 260 0 1 180
box -2 -2 2 2
use FILL  FILL_103
timestamp 1490995571
transform -1 0 256 0 1 90
box -8 -3 16 105
use FILL  FILL_104
timestamp 1490995571
transform -1 0 264 0 1 90
box -8 -3 16 105
use FILL  FILL_105
timestamp 1490995571
transform -1 0 272 0 1 90
box -8 -3 16 105
use FILL  FILL_106
timestamp 1490995571
transform -1 0 280 0 1 90
box -8 -3 16 105
use FILL  FILL_107
timestamp 1490995571
transform -1 0 288 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_188
timestamp 1490995571
transform 1 0 300 0 1 100
box -3 -3 3 3
use FILL  FILL_108
timestamp 1490995571
transform -1 0 296 0 1 90
box -8 -3 16 105
use FILL  FILL_109
timestamp 1490995571
transform -1 0 304 0 1 90
box -8 -3 16 105
use FILL  FILL_110
timestamp 1490995571
transform -1 0 312 0 1 90
box -8 -3 16 105
use FILL  FILL_111
timestamp 1490995571
transform -1 0 320 0 1 90
box -8 -3 16 105
use FILL  FILL_112
timestamp 1490995571
transform -1 0 328 0 1 90
box -8 -3 16 105
use FILL  FILL_113
timestamp 1490995571
transform -1 0 336 0 1 90
box -8 -3 16 105
use FILL  FILL_114
timestamp 1490995571
transform -1 0 344 0 1 90
box -8 -3 16 105
use FILL  FILL_115
timestamp 1490995571
transform -1 0 352 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_184
timestamp 1490995571
transform 1 0 364 0 1 180
box -3 -3 3 3
use FILL  FILL_116
timestamp 1490995571
transform -1 0 360 0 1 90
box -8 -3 16 105
use FILL  FILL_117
timestamp 1490995571
transform -1 0 368 0 1 90
box -8 -3 16 105
use FILL  FILL_118
timestamp 1490995571
transform -1 0 376 0 1 90
box -8 -3 16 105
use FILL  FILL_119
timestamp 1490995571
transform -1 0 384 0 1 90
box -8 -3 16 105
use FILL  FILL_120
timestamp 1490995571
transform -1 0 392 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_183
timestamp 1490995571
transform 1 0 428 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_185
timestamp 1490995571
transform 1 0 428 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_184
timestamp 1490995571
transform 1 0 412 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_185
timestamp 1490995571
transform 1 0 404 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_186
timestamp 1490995571
transform 1 0 404 0 1 110
box -3 -3 3 3
use FILL  FILL_121
timestamp 1490995571
transform -1 0 400 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_187
timestamp 1490995571
transform 1 0 428 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_189
timestamp 1490995571
transform 1 0 412 0 1 100
box -3 -3 3 3
use OR2X1  OR2X1_1
timestamp 1490995571
transform 1 0 400 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_186
timestamp 1490995571
transform 1 0 444 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_190
timestamp 1490995571
transform 1 0 444 0 1 180
box -3 -3 3 3
use FILL  FILL_122
timestamp 1490995571
transform -1 0 440 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_187
timestamp 1490995571
transform 1 0 452 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_188
timestamp 1490995571
transform 1 0 468 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_189
timestamp 1490995571
transform 1 0 460 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_191
timestamp 1490995571
transform 1 0 460 0 1 130
box -3 -3 3 3
use NAND3X1  NAND3X1_4
timestamp 1490995571
transform -1 0 472 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_190
timestamp 1490995571
transform 1 0 497 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_192
timestamp 1490995571
transform 1 0 497 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_199
timestamp 1490995571
transform 1 0 484 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_199
timestamp 1490995571
transform 1 0 484 0 1 110
box -3 -3 3 3
use FILL  FILL_123
timestamp 1490995571
transform -1 0 480 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_194
timestamp 1490995571
transform 1 0 508 0 1 139
box -2 -2 2 2
use $$M3_M2  $$M3_M2_193
timestamp 1490995571
transform 1 0 508 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_197
timestamp 1490995571
transform 1 0 500 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_196
timestamp 1490995571
transform 1 0 500 0 1 130
box -3 -3 3 3
use NOR2X1  NOR2X1_14
timestamp 1490995571
transform 1 0 480 0 1 90
box -8 -3 32 105
use FILL  FILL_124
timestamp 1490995571
transform -1 0 512 0 1 90
box -8 -3 16 105
use FILL  FILL_125
timestamp 1490995571
transform -1 0 520 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_195
timestamp 1490995571
transform 1 0 532 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_194
timestamp 1490995571
transform 1 0 532 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_200
timestamp 1490995571
transform 1 0 540 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_200
timestamp 1490995571
transform 1 0 540 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_15
timestamp 1490995571
transform -1 0 544 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_193
timestamp 1490995571
transform 1 0 580 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_196
timestamp 1490995571
transform 1 0 564 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_201
timestamp 1490995571
transform 1 0 556 0 1 110
box -3 -3 3 3
use FILL  FILL_126
timestamp 1490995571
transform -1 0 552 0 1 90
box -8 -3 16 105
use FILL  FILL_127
timestamp 1490995571
transform -1 0 560 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_195
timestamp 1490995571
transform 1 0 580 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_198
timestamp 1490995571
transform 1 0 572 0 1 134
box -2 -2 2 2
use $$M2_M1  $$M2_M1_191
timestamp 1490995571
transform 1 0 596 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_197
timestamp 1490995571
transform 1 0 588 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_198
timestamp 1490995571
transform 1 0 572 0 1 120
box -3 -3 3 3
use NAND3X1  NAND3X1_5
timestamp 1490995571
transform 1 0 560 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_192
timestamp 1490995571
transform 1 0 612 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_202
timestamp 1490995571
transform 1 0 604 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_201
timestamp 1490995571
transform 1 0 620 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_203
timestamp 1490995571
transform 1 0 620 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_202
timestamp 1490995571
transform 1 0 604 0 1 140
box -2 -2 2 2
use FILL  FILL_128
timestamp 1490995571
transform -1 0 600 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_204
timestamp 1490995571
transform 1 0 612 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_205
timestamp 1490995571
transform 1 0 628 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_203
timestamp 1490995571
transform 1 0 612 0 1 134
box -2 -2 2 2
use NAND3X1  NAND3X1_6
timestamp 1490995571
transform 1 0 600 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_204
timestamp 1490995571
transform 1 0 644 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_206
timestamp 1490995571
transform 1 0 644 0 1 150
box -3 -3 3 3
use FILL  FILL_129
timestamp 1490995571
transform -1 0 640 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_205
timestamp 1490995571
transform 1 0 660 0 1 130
box -2 -2 2 2
use $$M2_M1  $$M2_M1_206
timestamp 1490995571
transform 1 0 668 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_207
timestamp 1490995571
transform 1 0 668 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_208
timestamp 1490995571
transform 1 0 660 0 1 100
box -3 -3 3 3
use AND2X2  AND2X2_1
timestamp 1490995571
transform -1 0 672 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_209
timestamp 1490995571
transform 1 0 684 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_209
timestamp 1490995571
transform 1 0 684 0 1 127
box -2 -2 2 2
use FILL  FILL_130
timestamp 1490995571
transform -1 0 680 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_208
timestamp 1490995571
transform 1 0 692 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_210
timestamp 1490995571
transform 1 0 692 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_211
timestamp 1490995571
transform 1 0 700 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_210
timestamp 1490995571
transform 1 0 700 0 1 121
box -2 -2 2 2
use INVX2  INVX2_14
timestamp 1490995571
transform 1 0 680 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_207
timestamp 1490995571
transform 1 0 708 0 1 180
box -2 -2 2 2
use INVX2  INVX2_15
timestamp 1490995571
transform 1 0 696 0 1 90
box -9 -3 26 105
use FILL  FILL_131
timestamp 1490995571
transform -1 0 720 0 1 90
box -8 -3 16 105
use FILL  FILL_132
timestamp 1490995571
transform -1 0 728 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_212
timestamp 1490995571
transform 1 0 748 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_211
timestamp 1490995571
transform 1 0 740 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_213
timestamp 1490995571
transform 1 0 740 0 1 120
box -3 -3 3 3
use FILL  FILL_133
timestamp 1490995571
transform -1 0 736 0 1 90
box -8 -3 16 105
use FILL  FILL_134
timestamp 1490995571
transform -1 0 744 0 1 90
box -8 -3 16 105
use FILL  FILL_135
timestamp 1490995571
transform -1 0 752 0 1 90
box -8 -3 16 105
use FILL  FILL_136
timestamp 1490995571
transform -1 0 760 0 1 90
box -8 -3 16 105
use FILL  FILL_137
timestamp 1490995571
transform -1 0 768 0 1 90
box -8 -3 16 105
use INVX2  INVX2_16
timestamp 1490995571
transform -1 0 784 0 1 90
box -9 -3 26 105
use FILL  FILL_138
timestamp 1490995571
transform -1 0 792 0 1 90
box -8 -3 16 105
use FILL  FILL_139
timestamp 1490995571
transform -1 0 800 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_214
timestamp 1490995571
transform 1 0 812 0 1 150
box -3 -3 3 3
use FILL  FILL_140
timestamp 1490995571
transform -1 0 808 0 1 90
box -8 -3 16 105
use FILL  FILL_141
timestamp 1490995571
transform -1 0 816 0 1 90
box -8 -3 16 105
use FILL  FILL_142
timestamp 1490995571
transform -1 0 824 0 1 90
box -8 -3 16 105
use FILL  FILL_143
timestamp 1490995571
transform -1 0 832 0 1 90
box -8 -3 16 105
use FILL  FILL_144
timestamp 1490995571
transform -1 0 840 0 1 90
box -8 -3 16 105
use FILL  FILL_145
timestamp 1490995571
transform -1 0 848 0 1 90
box -8 -3 16 105
use FILL  FILL_146
timestamp 1490995571
transform -1 0 856 0 1 90
box -8 -3 16 105
use FILL  FILL_147
timestamp 1490995571
transform -1 0 864 0 1 90
box -8 -3 16 105
use FILL  FILL_148
timestamp 1490995571
transform -1 0 872 0 1 90
box -8 -3 16 105
use FILL  FILL_149
timestamp 1490995571
transform -1 0 880 0 1 90
box -8 -3 16 105
use FILL  FILL_150
timestamp 1490995571
transform -1 0 888 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_212
timestamp 1490995571
transform 1 0 900 0 1 130
box -2 -2 2 2
use FILL  FILL_151
timestamp 1490995571
transform -1 0 896 0 1 90
box -8 -3 16 105
use FILL  FILL_152
timestamp 1490995571
transform -1 0 904 0 1 90
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_9
timestamp 1490995571
transform 1 0 921 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1490995571
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1490995571
transform 1 0 921 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_215
timestamp 1490995571
transform 1 0 116 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_216
timestamp 1490995571
transform 1 0 884 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1490995571
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1490995571
transform 1 0 946 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 290 2 290 4 FreeSans 26 0 0 0 brnch
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 regdst
flabel metal3 2 170 2 170 4 FreeSans 26 0 0 0 regwrite
flabel metal3 2 520 2 520 4 FreeSans 26 0 0 0 iord
flabel metal3 2 400 2 400 4 FreeSans 26 0 0 0 pcwrite
flabel metal2 428 578 428 578 4 FreeSans 26 0 0 0 reset
flabel metal2 684 578 684 578 4 FreeSans 26 0 0 0 irwrite[3]
flabel metal2 44 578 44 578 4 FreeSans 26 0 0 0 memtoreg
flabel metal2 300 578 300 578 4 FreeSans 26 0 0 0 memwrite
flabel metal2 556 578 556 578 4 FreeSans 26 0 0 0 clk
flabel metal2 172 578 172 578 4 FreeSans 26 0 0 0 alusrca
flabel metal2 940 578 940 578 4 FreeSans 26 0 0 0 irwrite[1]
flabel metal2 812 578 812 578 4 FreeSans 26 0 0 0 irwrite[2]
flabel metal3 981 290 981 290 4 FreeSans 26 0 0 0 aluop[0]
flabel metal3 981 170 981 170 4 FreeSans 26 0 0 0 aluop[1]
flabel metal3 981 400 981 400 4 FreeSans 26 0 0 0 alusrcb[1]
flabel metal3 981 60 981 60 4 FreeSans 26 0 0 0 irwrite[0]
flabel metal3 981 520 981 520 4 FreeSans 26 0 0 0 alusrcb[0]
flabel metal2 172 1 172 1 4 FreeSans 26 0 0 0 pcsrc[0]
flabel metal2 428 1 428 1 4 FreeSans 26 0 0 0 op[4]
flabel metal2 684 1 684 1 4 FreeSans 26 0 0 0 op[2]
flabel metal2 300 1 300 1 4 FreeSans 26 0 0 0 op[5]
flabel metal2 812 1 812 1 4 FreeSans 26 0 0 0 op[1]
flabel metal2 556 1 556 1 4 FreeSans 26 0 0 0 op[3]
flabel metal2 940 1 940 1 4 FreeSans 26 0 0 0 op[0]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 pcsrc[1]
rlabel metal1 485 532 485 532 1 Vdd!
rlabel metal1 484 508 484 508 1 Gnd!
<< end >>
