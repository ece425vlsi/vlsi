magic
tech scmos
timestamp 1487096309
<< metal1 >>
rect -2 966 38 974
rect -2 876 38 884
rect 4 868 8 872
rect 44 868 48 872
<< m2contact >>
rect 0 868 4 872
rect 8 868 12 872
rect 40 868 44 872
rect 48 868 52 872
<< metal2 >>
rect 0 918 4 922
rect 8 872 12 922
rect 24 913 28 921
rect 32 918 36 922
rect 23 912 29 913
rect 23 908 24 912
rect 28 908 29 912
rect 23 907 29 908
rect 31 902 37 903
rect 31 898 32 902
rect 36 898 37 902
rect 31 897 37 898
rect 0 43 4 868
rect 32 50 36 897
rect 40 872 44 922
rect 56 903 60 921
rect 79 912 85 913
rect 79 908 80 912
rect 84 908 85 912
rect 79 907 85 908
rect 55 902 61 903
rect 55 898 56 902
rect 60 898 61 902
rect 55 897 61 898
rect 16 34 20 38
rect 24 34 28 38
rect 48 35 52 868
rect 80 57 84 907
rect 96 37 100 41
rect 72 33 76 37
<< m3contact >>
rect 24 908 28 912
rect 32 898 36 902
rect 80 908 84 912
rect 56 898 60 902
<< metal3 >>
rect 23 912 85 913
rect 23 908 24 912
rect 28 908 80 912
rect 84 908 85 912
rect 23 907 85 908
rect 31 902 61 903
rect 31 898 32 902
rect 36 898 56 902
rect 60 898 61 902
rect 31 897 61 898
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 0 0 1 880
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 32 0 1 880
box -6 -4 34 96
use mux4_dp_1x  mux4_dp_1x_0
timestamp 1484419186
transform 1 0 0 0 1 770
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_1
timestamp 1484419186
transform 1 0 0 0 1 660
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_2
timestamp 1484419186
transform 1 0 0 0 1 550
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_3
timestamp 1484419186
transform 1 0 0 0 1 440
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_4
timestamp 1484419186
transform 1 0 0 0 1 330
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_5
timestamp 1484419186
transform 1 0 0 0 1 220
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_6
timestamp 1484419186
transform 1 0 0 0 1 110
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_7
timestamp 1484419186
transform 1 0 0 0 1 0
box -6 -4 106 96
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 104 0 1 0
box -6 -4 130 866
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 232 0 1 0
box -6 -4 82 976
<< labels >>
rlabel metal2 0 918 4 922 1 s0
rlabel metal2 32 918 36 922 1 s1
rlabel metal2 16 34 20 38 1 d0_0_
rlabel metal2 24 34 28 38 1 d1_0_
rlabel metal2 72 33 76 37 1 d3_0_
rlabel metal2 96 37 100 41 1 y_0_
<< end >>
