magic
tech scmos
timestamp 1492530230
<< m2contact >>
rect -2 -2 2 2
<< end >>
