magic
tech scmos
timestamp 1488311656
<< m2contact >>
rect -2 -2 2 2
<< end >>
