magic
tech scmos
timestamp 1493737109
<< m2contact >>
rect -2 -2 2 2
<< end >>
