magic
tech scmos
timestamp 1493690834
<< metal2 >>
rect 1006 2222 1010 2459
rect 1013 2332 1017 2759
rect 1020 2442 1024 3059
rect 1027 2552 1031 3359
rect 1027 2547 1031 2548
rect 1020 2437 1024 2438
rect 1013 2327 1017 2328
rect 1006 2163 1010 2164
rect 1006 2112 1010 2159
rect 1020 2002 1024 2003
rect 1013 1892 1017 1893
rect 1006 1782 1010 1783
rect 1006 1050 1010 1778
rect 1013 1350 1017 1888
rect 1020 1863 1024 1998
rect 3350 1065 3354 1066
rect 1250 998 1254 1008
rect 1290 1007 1294 1008
rect 1394 1007 1398 1016
rect 1402 1007 1406 1025
rect 1550 1011 1554 1012
rect 1550 997 1554 1007
rect 1570 1006 1574 1034
rect 1578 1006 1582 1043
rect 1850 1020 1854 1021
rect 1850 998 1854 1016
rect 2122 1007 2126 1052
rect 2130 1007 2134 1061
rect 3050 1056 3054 1057
rect 2750 1047 2754 1048
rect 2150 1029 2154 1030
rect 2150 1000 2154 1025
rect 2150 998 2155 1000
rect 2450 998 2454 1034
rect 2750 998 2754 1043
rect 3050 998 3054 1052
rect 3350 1000 3354 1061
rect 3350 998 3355 1000
<< m3contact >>
rect 998 3359 1002 3363
rect 1027 3359 1031 3363
rect 998 3059 1002 3063
rect 1020 3059 1024 3063
rect 998 2759 1002 2763
rect 1013 2759 1017 2763
rect 998 2459 1002 2463
rect 1006 2459 1010 2463
rect 1027 2548 1031 2552
rect 1020 2438 1024 2442
rect 1013 2328 1017 2332
rect 1006 2218 1010 2222
rect 998 2159 1002 2163
rect 1006 2159 1010 2163
rect 1006 2108 1010 2112
rect 1020 1998 1024 2002
rect 1013 1888 1017 1892
rect 998 1859 1002 1863
rect 1006 1778 1010 1782
rect 998 1346 1002 1350
rect 1020 1859 1024 1863
rect 1013 1346 1017 1350
rect 2130 1061 2134 1065
rect 998 1046 1002 1050
rect 1006 1046 1010 1050
rect 2122 1052 2126 1056
rect 1578 1043 1582 1047
rect 1570 1034 1574 1038
rect 1402 1025 1406 1029
rect 1394 1016 1398 1020
rect 1250 1008 1254 1012
rect 1290 1008 1294 1012
rect 1386 1007 1390 1011
rect 1550 1007 1554 1011
rect 1850 1016 1854 1020
rect 3350 1061 3354 1065
rect 3050 1052 3054 1056
rect 2750 1043 2754 1047
rect 2450 1034 2454 1038
rect 2150 1025 2154 1029
<< metal3 >>
rect 997 3363 1032 3364
rect 997 3359 998 3363
rect 1002 3359 1027 3363
rect 1031 3359 1032 3363
rect 997 3358 1032 3359
rect 997 3063 1025 3064
rect 997 3059 998 3063
rect 1002 3059 1020 3063
rect 1024 3059 1025 3063
rect 997 3058 1025 3059
rect 997 2763 1018 2764
rect 997 2759 998 2763
rect 1002 2759 1013 2763
rect 1017 2759 1018 2763
rect 997 2758 1018 2759
rect 1007 2552 1186 2553
rect 1007 2548 1027 2552
rect 1031 2548 1186 2552
rect 1007 2547 1186 2548
rect 997 2463 1011 2464
rect 997 2459 998 2463
rect 1002 2459 1006 2463
rect 1010 2459 1011 2463
rect 997 2458 1011 2459
rect 1007 2442 1185 2443
rect 1007 2438 1020 2442
rect 1024 2438 1185 2442
rect 1007 2437 1185 2438
rect 1005 2332 1186 2333
rect 1005 2328 1013 2332
rect 1017 2328 1186 2332
rect 1005 2327 1186 2328
rect 1005 2222 1186 2223
rect 1005 2218 1006 2222
rect 1010 2218 1186 2222
rect 1005 2217 1186 2218
rect 997 2163 1011 2164
rect 997 2159 998 2163
rect 1002 2159 1006 2163
rect 1010 2159 1011 2163
rect 997 2158 1011 2159
rect 1005 2112 1186 2113
rect 1005 2108 1006 2112
rect 1010 2108 1186 2112
rect 1005 2107 1186 2108
rect 1007 2002 1185 2003
rect 1007 1998 1020 2002
rect 1024 1998 1185 2002
rect 1007 1997 1185 1998
rect 1007 1892 1185 1893
rect 1007 1888 1013 1892
rect 1017 1888 1185 1892
rect 1007 1887 1185 1888
rect 997 1863 1025 1864
rect 997 1859 998 1863
rect 1002 1859 1020 1863
rect 1024 1859 1025 1863
rect 997 1858 1025 1859
rect 1005 1782 1185 1783
rect 1005 1778 1006 1782
rect 1010 1778 1185 1782
rect 1005 1777 1185 1778
rect 997 1350 1018 1351
rect 997 1346 998 1350
rect 1002 1346 1013 1350
rect 1017 1346 1018 1350
rect 997 1345 1018 1346
rect 2129 1065 3355 1066
rect 2129 1061 2130 1065
rect 2134 1061 3350 1065
rect 3354 1061 3355 1065
rect 2129 1060 3355 1061
rect 2121 1056 3055 1057
rect 2121 1052 2122 1056
rect 2126 1052 3050 1056
rect 3054 1052 3055 1056
rect 2121 1051 3055 1052
rect 997 1050 1011 1051
rect 997 1046 998 1050
rect 1002 1046 1006 1050
rect 1010 1046 1011 1050
rect 997 1045 1011 1046
rect 1577 1047 2755 1048
rect 1577 1043 1578 1047
rect 1582 1043 2750 1047
rect 2754 1043 2755 1047
rect 1577 1042 2755 1043
rect 1569 1038 2455 1039
rect 1569 1034 1570 1038
rect 1574 1034 2450 1038
rect 2454 1034 2455 1038
rect 1569 1033 2455 1034
rect 1401 1029 2155 1030
rect 1401 1025 1402 1029
rect 1406 1025 2150 1029
rect 2154 1025 2155 1029
rect 1401 1024 2155 1025
rect 1393 1020 1855 1021
rect 1393 1016 1394 1020
rect 1398 1016 1850 1020
rect 1854 1016 1855 1020
rect 1393 1015 1855 1016
rect 1249 1012 1295 1013
rect 1249 1008 1250 1012
rect 1254 1008 1290 1012
rect 1294 1008 1295 1012
rect 1249 1007 1295 1008
rect 1385 1011 1555 1012
rect 1385 1007 1386 1011
rect 1390 1007 1550 1011
rect 1554 1007 1555 1011
rect 1385 1006 1555 1007
use alt_mips  alt_mips_0
timestamp 1493690834
transform 1 0 1115 0 1 1152
box 0 0 2876 1891
use PadFrame17  PadFrame17_0
timestamp 1491676833
transform 1 0 0 0 1 0
box 0 0 5000 5000
<< end >>
