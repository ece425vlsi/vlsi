magic
tech scmos
timestamp 1493737109
<< nwell >>
rect -8 48 64 105
<< ntransistor >>
rect 7 6 9 26
rect 16 6 18 26
rect 21 6 23 26
rect 33 6 35 26
rect 38 6 40 26
rect 47 6 49 26
<< ptransistor >>
rect 7 54 9 94
rect 16 54 18 94
rect 21 54 23 94
rect 33 54 35 94
rect 38 54 40 94
rect 47 54 49 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 21 16 26
rect 9 7 10 21
rect 14 7 16 21
rect 9 6 16 7
rect 18 6 21 26
rect 23 22 33 26
rect 23 8 26 22
rect 30 8 33 22
rect 23 6 33 8
rect 35 6 38 26
rect 40 21 47 26
rect 40 7 41 21
rect 45 7 47 21
rect 40 6 47 7
rect 49 25 54 26
rect 49 6 50 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 92 16 94
rect 9 63 10 92
rect 14 63 16 92
rect 9 54 16 63
rect 18 54 21 94
rect 23 93 33 94
rect 23 54 26 93
rect 30 54 33 93
rect 35 54 38 94
rect 40 92 47 94
rect 40 63 41 92
rect 45 63 47 92
rect 40 54 47 63
rect 49 93 54 94
rect 49 54 50 93
<< ndcontact >>
rect 2 6 6 25
rect 10 7 14 21
rect 26 8 30 22
rect 41 7 45 21
rect 50 6 54 25
<< pdcontact >>
rect 2 54 6 93
rect 10 63 14 92
rect 26 54 30 93
rect 41 63 45 92
rect 50 54 54 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
<< polysilicon >>
rect 7 94 9 96
rect 16 94 18 96
rect 21 94 23 96
rect 33 94 35 96
rect 38 94 40 96
rect 47 94 49 96
rect 7 37 9 54
rect 16 53 18 54
rect 15 51 18 53
rect 15 47 17 51
rect 7 26 9 33
rect 14 29 16 43
rect 21 39 23 54
rect 33 48 35 54
rect 38 53 40 54
rect 47 53 49 54
rect 38 51 49 53
rect 33 46 40 48
rect 38 37 40 46
rect 47 37 49 51
rect 24 35 32 37
rect 14 27 18 29
rect 16 26 18 27
rect 21 27 22 31
rect 30 29 32 35
rect 47 29 49 33
rect 30 27 35 29
rect 21 26 23 27
rect 33 26 35 27
rect 38 27 49 29
rect 38 26 40 27
rect 47 26 49 27
rect 7 4 9 6
rect 16 4 18 6
rect 21 4 23 6
rect 33 4 35 6
rect 38 4 40 6
rect 47 4 49 6
<< polycontact >>
rect 13 43 17 47
rect 6 33 10 37
rect 20 35 24 39
rect 22 27 26 31
rect 36 33 40 37
rect 46 33 50 37
<< metal1 >>
rect -2 102 58 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 58 102
rect -2 97 58 98
rect 11 94 15 97
rect 2 93 6 94
rect 10 92 15 94
rect 14 63 15 92
rect 10 61 15 63
rect 24 93 32 94
rect 6 54 11 57
rect 24 54 26 93
rect 30 54 32 93
rect 41 92 46 97
rect 45 63 46 92
rect 41 61 46 63
rect 50 93 54 94
rect 46 54 50 57
rect 27 47 30 54
rect 26 43 30 47
rect 2 33 6 37
rect 10 35 20 38
rect 27 37 30 43
rect 10 34 13 35
rect 27 34 32 37
rect 2 26 11 29
rect 2 25 6 26
rect 29 24 32 34
rect 50 33 54 37
rect 36 31 39 33
rect 46 26 54 29
rect 10 21 15 23
rect 14 7 15 21
rect 10 6 15 7
rect 24 22 32 24
rect 50 25 54 26
rect 24 8 26 22
rect 30 8 32 22
rect 24 6 32 8
rect 41 21 46 23
rect 45 7 46 21
rect 11 3 15 6
rect 41 3 46 7
rect -2 2 58 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 58 2
rect -2 -3 58 -2
<< m2contact >>
rect 11 54 15 58
rect 42 54 46 58
rect 17 44 21 48
rect 11 26 15 30
rect 18 27 22 31
rect 35 27 39 31
rect 42 26 46 30
<< metal2 >>
rect 11 30 14 54
rect 18 37 21 44
rect 43 37 46 54
rect 18 34 46 37
rect 15 27 18 30
rect 22 27 35 30
rect 43 30 46 34
<< labels >>
flabel metal1 28 45 28 45 4 FreeSans 26 0 0 0 Y
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 52 35 52 35 4 FreeSans 26 0 0 0 B
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
<< end >>
