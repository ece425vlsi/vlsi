magic
tech scmos
timestamp 1486490078
<< ntransistor >>
rect 7 7 9 23
rect 12 7 14 23
rect 17 7 19 23
<< ndiffusion >>
rect 2 22 7 23
rect 6 8 7 22
rect 2 7 7 8
rect 9 7 12 23
rect 14 7 17 23
rect 19 22 24 23
rect 19 8 20 22
rect 19 7 24 8
<< ndcontact >>
rect 2 8 6 22
rect 20 8 24 22
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< polysilicon >>
rect 7 23 9 31
rect 12 23 14 31
rect 17 23 19 31
rect 7 5 9 7
rect 12 5 14 7
rect 17 5 19 7
<< metal1 >>
rect 2 22 6 23
rect 2 4 6 8
rect 20 22 30 23
rect 24 19 30 22
rect 20 4 24 8
rect 0 2 32 4
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -4 32 -2
<< end >>
