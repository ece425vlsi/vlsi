magic
tech scmos
timestamp 1492562097
<< nwell >>
rect 280 44 290 100
<< psubstratepcontact >>
rect 278 2 282 6
rect 286 2 290 6
<< nsubstratencontact >>
rect 278 92 282 96
rect 286 92 290 96
<< polycontact >>
rect 326 142 330 146
rect 297 42 301 46
<< metal1 >>
rect 276 96 295 98
rect 276 92 278 96
rect 282 92 286 96
rect 290 92 295 96
rect 276 90 295 92
rect 275 6 295 8
rect 275 2 278 6
rect 282 2 286 6
rect 290 2 295 6
rect 275 0 295 2
<< m2contact >>
rect 608 220 612 224
rect 630 220 634 224
rect 652 220 656 224
rect 674 220 678 224
rect 696 220 700 224
rect 718 220 722 224
rect 740 220 744 224
rect 762 220 766 224
rect 593 196 597 200
rect 30 167 34 171
rect 110 167 114 171
rect 190 167 194 171
rect 270 167 274 171
rect 350 167 354 171
rect 430 167 434 171
rect 510 167 514 171
rect 593 168 597 172
rect 326 142 330 146
rect 406 142 410 146
rect 486 142 490 146
rect 593 140 597 144
rect 593 112 597 116
rect 593 84 597 88
rect 593 56 597 60
rect 230 50 234 54
rect 304 51 308 55
rect 198 42 202 46
rect 270 42 274 46
rect 296 42 297 46
rect 297 42 300 46
rect 593 28 597 32
rect 593 0 597 4
rect 619 0 623 4
rect 641 0 645 4
rect 663 0 667 4
rect 685 0 689 4
rect 707 0 711 4
rect 729 0 733 4
rect 751 0 755 4
<< metal2 >>
rect 6 155 10 238
rect 14 159 18 229
rect 22 159 26 214
rect 6 -59 10 46
rect 14 38 18 151
rect 38 127 42 155
rect 31 16 35 69
rect 38 -50 42 46
rect 45 32 49 104
rect 54 34 58 301
rect 70 108 74 163
rect 94 159 98 229
rect 102 159 106 214
rect 134 155 138 301
rect 94 136 98 151
rect 63 16 67 69
rect 70 -41 74 46
rect 86 34 90 132
rect 118 127 122 155
rect 95 16 99 69
rect 102 -32 106 46
rect 118 34 122 57
rect 127 16 131 69
rect 134 -23 138 46
rect 142 38 146 132
rect 150 78 154 163
rect 174 159 178 229
rect 182 159 186 214
rect 198 127 202 155
rect 142 34 154 38
rect 159 16 163 69
rect 166 -14 170 46
rect 182 34 186 114
rect 191 16 195 69
rect 198 -5 202 42
rect 206 38 210 105
rect 214 61 218 301
rect 246 242 250 301
rect 230 87 234 163
rect 246 155 250 238
rect 254 159 258 229
rect 223 46 227 69
rect 238 63 242 151
rect 230 54 234 59
rect 206 34 218 38
rect 223 16 227 42
rect 238 46 242 54
rect 262 48 266 214
rect 278 127 282 155
rect 294 136 298 301
rect 326 242 330 243
rect 310 96 314 163
rect 318 162 322 163
rect 326 162 330 238
rect 318 109 322 158
rect 334 65 338 229
rect 342 159 346 214
rect 344 127 348 129
rect 358 127 362 155
rect 296 46 300 61
rect 344 46 348 123
rect 374 118 378 301
rect 454 242 458 301
rect 390 105 394 163
rect 414 159 418 229
rect 422 218 426 219
rect 422 159 426 214
rect 454 167 458 238
rect 470 159 474 179
rect 494 159 498 229
rect 534 218 538 301
rect 502 159 506 214
rect 534 167 538 214
rect 550 200 555 201
rect 554 196 555 200
rect 550 159 555 196
rect 561 178 565 301
rect 585 233 589 300
rect 600 223 604 300
rect 608 224 612 291
rect 622 223 626 300
rect 630 224 634 282
rect 644 223 648 300
rect 652 224 656 273
rect 666 223 670 300
rect 674 224 678 264
rect 688 223 692 300
rect 696 224 700 255
rect 710 223 714 300
rect 718 224 722 246
rect 732 223 736 300
rect 740 224 744 237
rect 754 223 758 300
rect 762 224 766 228
rect 608 194 609 198
rect 613 194 765 198
rect 561 174 572 178
rect 561 167 562 171
rect 568 163 572 174
rect 579 172 583 179
rect 561 159 572 163
rect 438 127 442 155
rect 518 127 522 155
rect 561 146 565 159
rect 572 105 576 140
rect 581 96 585 112
rect 559 60 563 74
rect 238 16 242 42
rect 280 4 284 42
rect 776 47 780 228
rect 296 16 300 42
rect 619 -5 623 0
rect 641 -14 645 0
rect 663 -23 667 0
rect 685 -32 689 0
rect 707 -41 711 0
rect 729 -50 733 0
rect 751 -59 755 0
rect 783 -43 787 237
rect 790 -23 794 246
rect 797 -3 801 255
rect 804 27 808 264
rect 811 67 815 273
rect 818 97 822 282
rect 825 127 829 291
rect 853 198 857 199
rect 853 157 857 194
rect 860 177 864 300
rect 867 217 871 300
rect 874 197 878 300
<< m3contact >>
rect 6 238 10 242
rect 14 229 18 233
rect 22 214 26 218
rect 6 151 10 155
rect 14 151 18 155
rect 6 142 10 146
rect 38 123 42 127
rect 45 104 49 108
rect 14 34 18 38
rect 22 34 26 38
rect 31 12 35 16
rect 94 229 98 233
rect 102 214 106 218
rect 174 229 178 233
rect 94 151 98 155
rect 86 142 90 146
rect 70 104 74 108
rect 86 132 90 136
rect 94 132 98 136
rect 45 28 49 32
rect 63 12 67 16
rect 134 151 138 155
rect 118 123 122 127
rect 142 132 146 136
rect 118 57 122 61
rect 95 12 99 16
rect 127 12 131 16
rect 182 214 186 218
rect 166 142 170 146
rect 198 123 202 127
rect 150 74 154 78
rect 182 114 186 118
rect 159 12 163 16
rect 206 105 210 109
rect 191 12 195 16
rect 246 238 250 242
rect 254 229 258 233
rect 262 214 266 218
rect 230 83 234 87
rect 238 151 242 155
rect 246 151 250 155
rect 214 57 218 61
rect 246 142 250 146
rect 230 59 234 63
rect 238 59 242 63
rect 254 59 258 63
rect 223 42 227 46
rect 223 12 227 16
rect 326 238 330 242
rect 294 132 298 136
rect 278 123 282 127
rect 318 158 322 162
rect 326 158 330 162
rect 334 229 338 233
rect 326 142 330 146
rect 318 105 322 109
rect 310 92 314 96
rect 342 214 346 218
rect 296 61 300 65
rect 334 61 338 65
rect 344 123 348 127
rect 358 123 362 127
rect 304 51 308 55
rect 454 238 458 242
rect 414 229 418 233
rect 374 114 378 118
rect 422 214 426 218
rect 494 229 498 233
rect 470 179 474 183
rect 502 214 506 218
rect 534 214 538 218
rect 550 196 554 200
rect 585 229 589 233
rect 600 219 604 223
rect 608 291 612 295
rect 622 219 626 223
rect 630 282 634 286
rect 644 219 648 223
rect 652 273 656 277
rect 666 219 670 223
rect 674 264 678 268
rect 688 219 692 223
rect 696 255 700 259
rect 710 219 714 223
rect 718 246 722 250
rect 732 219 736 223
rect 740 237 744 241
rect 825 291 829 295
rect 818 282 822 286
rect 811 273 815 277
rect 804 264 808 268
rect 797 255 801 259
rect 790 246 794 250
rect 783 237 787 241
rect 754 219 758 223
rect 762 228 766 232
rect 776 228 780 232
rect 600 212 604 216
rect 593 196 597 200
rect 609 194 613 198
rect 765 194 769 198
rect 622 184 626 188
rect 579 179 583 183
rect 579 168 583 172
rect 593 168 597 172
rect 406 142 410 146
rect 486 142 490 146
rect 438 123 442 127
rect 644 156 648 160
rect 561 142 565 146
rect 518 123 522 127
rect 572 140 576 144
rect 593 140 597 144
rect 390 101 394 105
rect 666 128 670 132
rect 572 101 576 105
rect 581 112 585 116
rect 593 112 597 116
rect 688 100 692 104
rect 581 92 585 96
rect 593 84 597 88
rect 559 74 563 78
rect 710 72 714 76
rect 559 56 563 60
rect 593 56 597 60
rect 238 42 242 46
rect 270 42 274 46
rect 280 42 284 46
rect 238 12 242 16
rect 304 42 308 46
rect 344 42 348 46
rect 732 44 736 48
rect 776 43 780 47
rect 593 28 597 32
rect 754 16 758 20
rect 296 12 300 16
rect 280 0 284 4
rect 593 0 597 4
rect 198 -9 202 -5
rect 619 -9 623 -5
rect 166 -18 170 -14
rect 641 -18 645 -14
rect 134 -27 138 -23
rect 663 -27 667 -23
rect 102 -36 106 -32
rect 685 -36 689 -32
rect 70 -45 74 -41
rect 707 -45 711 -41
rect 38 -54 42 -50
rect 729 -54 733 -50
rect 6 -63 10 -59
rect 853 194 857 198
rect 867 213 871 217
rect 874 193 878 197
rect 860 173 864 177
rect 853 153 857 157
rect 825 123 829 127
rect 818 93 822 97
rect 811 63 815 67
rect 804 23 808 27
rect 797 -7 801 -3
rect 790 -27 794 -23
rect 783 -47 787 -43
rect 751 -63 755 -59
<< metal3 >>
rect 607 295 830 296
rect 607 291 608 295
rect 612 291 825 295
rect 829 291 830 295
rect 607 290 830 291
rect 629 286 823 287
rect 629 282 630 286
rect 634 282 818 286
rect 822 282 823 286
rect 629 281 823 282
rect 651 277 816 278
rect 651 273 652 277
rect 656 273 811 277
rect 815 273 816 277
rect 651 272 816 273
rect 673 268 809 269
rect 673 264 674 268
rect 678 264 804 268
rect 808 264 809 268
rect 673 263 809 264
rect 695 259 802 260
rect 695 255 696 259
rect 700 255 797 259
rect 801 255 802 259
rect 695 254 802 255
rect 717 250 795 251
rect 717 246 718 250
rect 722 246 790 250
rect 794 246 795 250
rect 717 245 795 246
rect 5 242 251 243
rect 5 238 6 242
rect 10 238 246 242
rect 250 238 251 242
rect 5 237 251 238
rect 325 242 459 243
rect 325 238 326 242
rect 330 238 454 242
rect 458 238 459 242
rect 325 237 459 238
rect 739 241 788 242
rect 739 237 740 241
rect 744 237 783 241
rect 787 237 788 241
rect 739 236 788 237
rect 13 233 614 234
rect 13 229 14 233
rect 18 229 94 233
rect 98 229 174 233
rect 178 229 254 233
rect 258 229 334 233
rect 338 229 414 233
rect 418 229 494 233
rect 498 229 585 233
rect 589 229 614 233
rect 13 228 614 229
rect 599 223 605 224
rect 599 219 600 223
rect 604 219 605 223
rect 21 218 539 219
rect 21 214 22 218
rect 26 214 102 218
rect 106 214 182 218
rect 186 214 262 218
rect 266 214 342 218
rect 346 214 422 218
rect 426 214 502 218
rect 506 214 534 218
rect 538 214 539 218
rect 21 213 539 214
rect 599 216 605 219
rect 599 212 600 216
rect 604 212 605 216
rect 599 211 605 212
rect 549 200 598 201
rect 549 196 550 200
rect 554 196 593 200
rect 597 196 598 200
rect 549 195 598 196
rect 608 198 614 228
rect 761 232 781 233
rect 761 228 762 232
rect 766 228 776 232
rect 780 228 781 232
rect 761 227 781 228
rect 608 194 609 198
rect 613 194 614 198
rect 608 193 614 194
rect 621 223 627 224
rect 621 219 622 223
rect 626 219 627 223
rect 621 188 627 219
rect 621 184 622 188
rect 626 184 627 188
rect 469 183 584 184
rect 621 183 627 184
rect 643 223 649 224
rect 643 219 644 223
rect 648 219 649 223
rect 469 179 470 183
rect 474 179 579 183
rect 583 179 584 183
rect 469 178 584 179
rect 578 172 598 173
rect 578 168 579 172
rect 583 168 593 172
rect 597 168 598 172
rect 578 167 598 168
rect 317 162 331 163
rect 317 158 318 162
rect 322 158 326 162
rect 330 158 331 162
rect 317 157 331 158
rect 643 160 649 219
rect 643 156 644 160
rect 648 156 649 160
rect 5 155 19 156
rect 5 151 6 155
rect 10 151 14 155
rect 18 151 19 155
rect 5 150 19 151
rect 93 155 139 156
rect 93 151 94 155
rect 98 151 134 155
rect 138 151 139 155
rect 93 150 139 151
rect 237 155 251 156
rect 643 155 649 156
rect 665 223 671 224
rect 665 219 666 223
rect 670 219 671 223
rect 237 151 238 155
rect 242 151 246 155
rect 250 151 251 155
rect 237 150 251 151
rect 5 146 566 147
rect 5 142 6 146
rect 10 142 86 146
rect 90 142 166 146
rect 170 142 246 146
rect 250 142 326 146
rect 330 142 406 146
rect 410 142 486 146
rect 490 142 561 146
rect 565 142 566 146
rect 5 141 566 142
rect 571 144 598 145
rect 571 140 572 144
rect 576 140 593 144
rect 597 140 598 144
rect 571 139 598 140
rect 85 136 99 137
rect 85 132 86 136
rect 90 132 94 136
rect 98 132 99 136
rect 85 131 99 132
rect 141 136 299 137
rect 141 132 142 136
rect 146 132 294 136
rect 298 132 299 136
rect 141 131 299 132
rect 665 132 671 219
rect 665 128 666 132
rect 670 128 671 132
rect 35 127 523 128
rect 665 127 671 128
rect 687 223 693 224
rect 687 219 688 223
rect 692 219 693 223
rect 35 123 38 127
rect 42 123 118 127
rect 122 123 198 127
rect 202 123 278 127
rect 282 123 344 127
rect 348 123 358 127
rect 362 123 438 127
rect 442 123 518 127
rect 522 123 523 127
rect 35 122 523 123
rect 181 118 379 119
rect 181 114 182 118
rect 186 114 374 118
rect 378 114 379 118
rect 181 113 379 114
rect 580 116 598 117
rect 580 112 581 116
rect 585 112 593 116
rect 597 112 598 116
rect 580 111 598 112
rect 205 109 323 110
rect 44 108 75 109
rect 44 104 45 108
rect 49 104 70 108
rect 74 104 75 108
rect 205 105 206 109
rect 210 105 318 109
rect 322 105 323 109
rect 205 104 323 105
rect 389 105 577 106
rect 44 103 75 104
rect 389 101 390 105
rect 394 101 572 105
rect 576 101 577 105
rect 389 100 577 101
rect 687 104 693 219
rect 687 100 688 104
rect 692 100 693 104
rect 687 99 693 100
rect 709 223 715 224
rect 709 219 710 223
rect 714 219 715 223
rect 309 96 586 97
rect 309 92 310 96
rect 314 92 581 96
rect 585 92 586 96
rect 309 91 586 92
rect 592 88 598 89
rect 229 87 593 88
rect 229 83 230 87
rect 234 84 593 87
rect 597 84 598 88
rect 234 83 598 84
rect 229 82 598 83
rect 149 78 564 79
rect 149 74 150 78
rect 154 74 559 78
rect 563 74 564 78
rect 149 73 564 74
rect 709 76 715 219
rect 709 72 710 76
rect 714 72 715 76
rect 709 71 715 72
rect 731 223 737 224
rect 731 219 732 223
rect 736 219 737 223
rect 295 65 339 66
rect 229 63 243 64
rect 117 61 219 62
rect 117 57 118 61
rect 122 57 214 61
rect 218 57 219 61
rect 229 59 230 63
rect 234 59 238 63
rect 242 59 243 63
rect 229 58 243 59
rect 253 63 285 64
rect 253 59 254 63
rect 258 59 285 63
rect 295 61 296 65
rect 300 61 334 65
rect 338 61 339 65
rect 295 60 339 61
rect 558 60 598 61
rect 253 58 285 59
rect 117 56 219 57
rect 279 56 285 58
rect 558 56 559 60
rect 563 56 593 60
rect 597 56 598 60
rect 279 55 309 56
rect 558 55 598 56
rect 279 51 304 55
rect 308 51 309 55
rect 279 50 309 51
rect 731 48 737 219
rect 222 46 243 47
rect 222 42 223 46
rect 227 42 238 46
rect 242 42 243 46
rect 222 41 243 42
rect 269 46 285 47
rect 269 42 270 46
rect 274 42 280 46
rect 284 42 285 46
rect 269 41 285 42
rect 303 46 349 47
rect 303 42 304 46
rect 308 42 344 46
rect 348 42 349 46
rect 731 44 732 48
rect 736 44 737 48
rect 731 43 737 44
rect 753 223 759 224
rect 753 219 754 223
rect 758 219 759 223
rect 303 41 349 42
rect 13 38 27 39
rect 13 34 14 38
rect 18 34 22 38
rect 26 34 27 38
rect 13 33 27 34
rect 44 32 598 33
rect 44 28 45 32
rect 49 28 593 32
rect 597 28 598 32
rect 44 27 598 28
rect 753 20 759 219
rect 866 217 879 218
rect 866 213 867 217
rect 871 213 879 217
rect 866 212 879 213
rect 764 198 858 199
rect 764 194 765 198
rect 769 194 853 198
rect 857 194 858 198
rect 764 193 858 194
rect 873 197 879 198
rect 873 193 874 197
rect 878 193 879 197
rect 873 192 879 193
rect 859 177 879 178
rect 859 173 860 177
rect 864 173 879 177
rect 859 172 879 173
rect 852 157 879 158
rect 852 153 853 157
rect 857 153 879 157
rect 852 152 879 153
rect 824 127 881 128
rect 824 123 825 127
rect 829 123 881 127
rect 824 122 830 123
rect 817 97 879 98
rect 817 93 818 97
rect 822 93 879 97
rect 817 92 823 93
rect 810 67 876 68
rect 810 63 811 67
rect 815 63 876 67
rect 810 62 816 63
rect 775 47 875 48
rect 775 43 776 47
rect 780 43 875 47
rect 775 42 781 43
rect 803 27 876 28
rect 803 23 804 27
rect 808 23 876 27
rect 803 22 809 23
rect 30 16 228 17
rect 30 12 31 16
rect 35 12 63 16
rect 67 12 95 16
rect 99 12 127 16
rect 131 12 159 16
rect 163 12 191 16
rect 195 12 223 16
rect 227 12 228 16
rect 30 11 228 12
rect 237 16 301 17
rect 237 12 238 16
rect 242 12 296 16
rect 300 12 301 16
rect 753 16 754 20
rect 758 16 759 20
rect 753 15 759 16
rect 237 11 301 12
rect 279 4 598 5
rect 279 0 280 4
rect 284 0 593 4
rect 597 0 598 4
rect 279 -1 598 0
rect 796 -3 874 -2
rect 197 -5 624 -4
rect 197 -9 198 -5
rect 202 -9 619 -5
rect 623 -9 624 -5
rect 796 -7 797 -3
rect 801 -7 874 -3
rect 796 -8 802 -7
rect 197 -10 624 -9
rect 165 -14 646 -13
rect 165 -18 166 -14
rect 170 -18 641 -14
rect 645 -18 646 -14
rect 165 -19 646 -18
rect 133 -23 668 -22
rect 133 -27 134 -23
rect 138 -27 663 -23
rect 667 -27 668 -23
rect 133 -28 668 -27
rect 789 -23 874 -22
rect 789 -27 790 -23
rect 794 -27 874 -23
rect 789 -28 795 -27
rect 101 -32 690 -31
rect 101 -36 102 -32
rect 106 -36 685 -32
rect 689 -36 690 -32
rect 101 -37 690 -36
rect 69 -41 712 -40
rect 69 -45 70 -41
rect 74 -45 707 -41
rect 711 -45 712 -41
rect 69 -46 712 -45
rect 782 -43 875 -42
rect 782 -47 783 -43
rect 787 -47 875 -43
rect 782 -48 788 -47
rect 37 -50 734 -49
rect 37 -54 38 -50
rect 42 -54 729 -50
rect 733 -54 734 -50
rect 37 -55 734 -54
rect 5 -59 756 -58
rect 5 -63 6 -59
rect 10 -63 751 -59
rect 755 -63 756 -59
rect 5 -64 756 -63
use inv_1x  inv_1x_0
timestamp 1492544053
transform 1 0 296 0 1 4
box -6 -4 18 96
use source_gen_7_0  source_gen_7_0_0
timestamp 1492561529
transform 1 0 0 0 1 0
box 0 0 773 224
use three_eight_decoder  three_eight_decoder_0
timestamp 1492530230
transform 1 0 873 0 1 -104
box 0 40 666 340
<< labels >>
rlabel metal2 536 299 536 299 5 a7
rlabel metal2 456 299 456 299 5 a6
rlabel metal2 376 299 376 299 5 a5
rlabel metal2 296 299 296 299 5 a4
rlabel metal2 216 299 216 299 5 a3
rlabel metal2 136 299 136 299 5 a2
rlabel metal2 56 299 56 299 5 a1
rlabel metal2 587 297 587 297 5 right
rlabel metal2 563 299 563 299 5 arith
rlabel metal2 248 299 248 299 5 a0
rlabel metal2 602 298 602 298 5 y7
rlabel metal2 624 298 624 298 5 y6
rlabel metal2 646 298 646 298 5 y5
rlabel metal2 668 298 668 298 5 y4
rlabel metal2 690 298 690 298 5 y3
rlabel metal2 712 298 712 298 5 y2
rlabel metal2 734 298 734 298 5 y1
rlabel metal2 756 298 756 298 5 y0
rlabel metal2 869 298 869 298 5 k1
rlabel metal2 876 298 876 298 5 k0
rlabel metal2 862 298 862 298 5 k2
rlabel space 1021 229 1021 229 1 Vdd!
rlabel space 1021 204 1021 204 1 Gnd!
rlabel space 76 206 76 206 1 Vdd!
rlabel space 76 116 76 116 1 Gnd!
rlabel space 76 94 76 94 1 Vdd!
rlabel space 76 4 76 4 1 Gnd!
rlabel metal3 863 125 863 125 1 s7
rlabel metal3 859 95 859 95 1 s6
rlabel metal3 858 65 858 65 1 s5
rlabel metal3 857 45 857 45 1 s0
rlabel metal3 861 26 861 26 1 s4
rlabel metal3 856 -5 856 -5 1 s3
rlabel metal3 857 -25 857 -25 1 s2
rlabel metal3 857 -45 857 -45 1 s1
rlabel metal3 743 -61 743 -61 1 z0
rlabel metal3 722 -53 722 -53 1 z1
rlabel metal3 701 -44 701 -44 1 z2
rlabel metal3 676 -34 676 -34 1 z3
rlabel metal3 653 -25 653 -25 1 z4
rlabel metal3 632 -17 632 -17 1 z5
rlabel metal3 605 -8 605 -8 1 z6
rlabel metal3 585 2 585 2 1 z7
rlabel metal3 584 31 584 31 1 z8
rlabel metal3 584 58 584 58 1 z9
rlabel metal3 583 84 583 84 1 z10
rlabel metal3 575 93 575 93 1 z11
rlabel metal3 564 103 564 103 1 z12
rlabel metal3 588 171 588 171 1 z13
rlabel metal3 589 199 589 199 1 z14
rlabel metal3 319 43 319 43 1 rightb
rlabel metal3 276 42 276 42 1 zout
rlabel metal2 264 54 264 54 1 a7in
rlabel metal2 231 56 231 56 1 a0in
<< end >>
