magic
tech scmos
timestamp 1490995571
<< m2contact >>
rect -7 -2 7 2
<< end >>
