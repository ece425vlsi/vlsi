magic
tech scmos
timestamp 1493740799
<< metal2 >>
rect 564 1941 568 1942
rect 380 1932 384 1933
rect 364 1923 368 1924
rect 356 1914 360 1915
rect 348 1905 352 1906
rect 340 1896 344 1897
rect 332 1887 336 1888
rect 324 1878 328 1879
rect 196 1869 200 1870
rect 140 1860 144 1861
rect 196 1859 200 1865
rect 324 1856 328 1874
rect 332 1858 336 1883
rect 340 1856 344 1892
rect 348 1856 352 1901
rect 356 1855 360 1910
rect 364 1856 368 1919
rect 380 1853 384 1928
rect 564 1854 568 1937
rect 581 1860 585 1952
rect 605 1869 609 1952
rect 637 1878 641 1952
rect 669 1887 673 1952
rect 709 1896 713 1952
rect 741 1905 745 1952
rect 773 1914 777 1952
rect 805 1923 809 1952
rect 837 1932 841 1952
rect 869 1941 873 1952
rect 869 1936 873 1937
rect 837 1927 841 1928
rect 852 1932 856 1933
rect 805 1918 809 1919
rect 836 1923 840 1924
rect 773 1909 777 1910
rect 741 1900 745 1901
rect 709 1891 713 1892
rect 724 1896 728 1897
rect 669 1882 673 1883
rect 637 1873 641 1874
rect 605 1864 609 1865
rect 724 1859 728 1892
rect 836 1856 840 1919
rect 852 1858 856 1928
rect 860 1914 864 1915
rect 860 1859 864 1910
rect 868 1905 872 1906
rect 868 1856 872 1901
rect 909 1896 913 1952
rect 941 1923 945 1952
rect 973 1932 977 1952
rect 973 1927 977 1928
rect 941 1918 945 1919
rect 1005 1914 1009 1952
rect 1005 1909 1009 1910
rect 1037 1905 1041 1952
rect 1037 1900 1041 1901
rect 909 1891 913 1892
rect 876 1887 880 1888
rect 876 1859 880 1883
rect 1069 1887 1073 1952
rect 1069 1882 1073 1883
rect 884 1878 888 1879
rect 884 1859 888 1874
rect 1109 1878 1113 1952
rect 1109 1873 1113 1874
rect 892 1869 896 1870
rect 892 1859 896 1865
rect 1141 1869 1145 1952
rect 1141 1864 1145 1865
<< m3contact >>
rect 564 1937 568 1941
rect 380 1928 384 1932
rect 364 1919 368 1923
rect 356 1910 360 1914
rect 348 1901 352 1905
rect 340 1892 344 1896
rect 332 1883 336 1887
rect 324 1874 328 1878
rect 196 1865 200 1869
rect 140 1856 144 1860
rect 869 1937 873 1941
rect 837 1928 841 1932
rect 852 1928 856 1932
rect 805 1919 809 1923
rect 836 1919 840 1923
rect 773 1910 777 1914
rect 741 1901 745 1905
rect 709 1892 713 1896
rect 724 1892 728 1896
rect 669 1883 673 1887
rect 637 1874 641 1878
rect 605 1865 609 1869
rect 581 1856 585 1860
rect 860 1910 864 1914
rect 868 1901 872 1905
rect 973 1928 977 1932
rect 941 1919 945 1923
rect 1005 1910 1009 1914
rect 1037 1901 1041 1905
rect 909 1892 913 1896
rect 876 1883 880 1887
rect 1069 1883 1073 1887
rect 884 1874 888 1878
rect 1109 1874 1113 1878
rect 892 1865 896 1869
rect 1141 1865 1145 1869
<< metal3 >>
rect 563 1941 874 1942
rect 563 1937 564 1941
rect 568 1937 869 1941
rect 873 1937 874 1941
rect 563 1936 874 1937
rect 379 1932 842 1933
rect 379 1928 380 1932
rect 384 1928 837 1932
rect 841 1928 842 1932
rect 379 1927 842 1928
rect 851 1932 978 1933
rect 851 1928 852 1932
rect 856 1928 973 1932
rect 977 1928 978 1932
rect 851 1927 978 1928
rect 363 1923 810 1924
rect 363 1919 364 1923
rect 368 1919 805 1923
rect 809 1919 810 1923
rect 363 1918 810 1919
rect 835 1923 946 1924
rect 835 1919 836 1923
rect 840 1919 941 1923
rect 945 1919 946 1923
rect 835 1918 946 1919
rect 355 1914 778 1915
rect 355 1910 356 1914
rect 360 1910 773 1914
rect 777 1910 778 1914
rect 355 1909 778 1910
rect 859 1914 1010 1915
rect 859 1910 860 1914
rect 864 1910 1005 1914
rect 1009 1910 1010 1914
rect 859 1909 1010 1910
rect 347 1905 746 1906
rect 347 1901 348 1905
rect 352 1901 741 1905
rect 745 1901 746 1905
rect 347 1900 746 1901
rect 867 1905 1042 1906
rect 867 1901 868 1905
rect 872 1901 1037 1905
rect 1041 1901 1042 1905
rect 867 1900 1042 1901
rect 339 1896 714 1897
rect 339 1892 340 1896
rect 344 1892 709 1896
rect 713 1892 714 1896
rect 339 1891 714 1892
rect 723 1896 914 1897
rect 723 1892 724 1896
rect 728 1892 909 1896
rect 913 1892 914 1896
rect 723 1891 914 1892
rect 331 1887 674 1888
rect 331 1883 332 1887
rect 336 1883 669 1887
rect 673 1883 674 1887
rect 331 1882 674 1883
rect 875 1887 1074 1888
rect 875 1883 876 1887
rect 880 1883 1069 1887
rect 1073 1883 1074 1887
rect 875 1882 1074 1883
rect 323 1878 642 1879
rect 323 1874 324 1878
rect 328 1874 637 1878
rect 641 1874 642 1878
rect 323 1873 642 1874
rect 883 1878 1114 1879
rect 883 1874 884 1878
rect 888 1874 1109 1878
rect 1113 1874 1114 1878
rect 883 1873 1114 1874
rect 195 1869 610 1870
rect 195 1865 196 1869
rect 200 1865 605 1869
rect 609 1865 610 1869
rect 195 1864 610 1865
rect 891 1869 1146 1870
rect 891 1865 892 1869
rect 896 1865 1141 1869
rect 1145 1865 1146 1869
rect 891 1864 1146 1865
rect 139 1860 586 1861
rect 139 1856 140 1860
rect 144 1856 581 1860
rect 585 1856 586 1860
rect 139 1855 586 1856
use alt_controller  alt_controller_0
timestamp 1493737109
transform 1 0 540 0 1 1952
box 0 0 2082 380
use datapath  datapath_0
timestamp 1493739066
transform 1 0 140 0 1 548
box -140 -548 2736 1343
<< end >>
