magic
tech scmos
timestamp 1493691729
<< metal1 >>
rect -140 1302 2664 1304
rect -76 1298 2600 1302
rect -140 1296 2664 1298
rect 817 1248 827 1252
rect -68 1212 2736 1214
rect -4 1208 2672 1212
rect -68 1206 2736 1208
rect 820 1198 856 1202
rect 876 1198 888 1202
rect -140 1192 2664 1194
rect -76 1188 2600 1192
rect -140 1186 2664 1188
rect -68 1102 2736 1104
rect -4 1098 2672 1102
rect -68 1096 2736 1098
rect 820 1088 872 1092
rect -140 1082 2664 1084
rect -76 1078 2600 1082
rect -140 1076 2664 1078
rect -68 992 2736 994
rect -4 988 2672 992
rect -68 986 2736 988
rect 2451 974 2455 976
rect 2527 974 2531 976
rect -140 972 2664 974
rect -76 968 2600 972
rect -140 966 2461 968
rect 2473 966 2477 968
rect 2497 966 2501 968
rect 2513 966 2517 968
rect 2528 966 2664 968
rect -68 882 2736 884
rect -4 878 2672 882
rect -68 876 2736 878
rect -140 862 2231 864
rect -76 858 2231 862
rect -140 856 2231 858
rect 2479 862 2664 864
rect 2479 858 2600 862
rect 2479 856 2664 858
rect 856 816 875 820
rect 177 812 184 816
rect 361 812 368 816
rect 856 813 860 816
rect 1808 815 1812 819
rect 1801 811 1812 815
rect 2032 812 2067 816
rect 2032 808 2036 812
rect -68 772 2231 774
rect -4 771 2231 772
rect -4 768 1624 771
rect -68 767 1624 768
rect 1628 767 2231 771
rect -68 766 2231 767
rect 2479 772 2736 774
rect 2479 768 2672 772
rect 2479 766 2736 768
rect 1668 757 1672 761
rect -140 752 2199 754
rect -76 748 2199 752
rect -140 746 2199 748
rect 2479 752 2664 754
rect 2479 748 2600 752
rect 2479 746 2664 748
rect 856 706 875 710
rect 177 702 192 706
rect 361 702 376 706
rect 856 703 860 706
rect 1808 705 1812 709
rect 1801 701 1812 705
rect 2032 702 2067 706
rect 2032 698 2036 702
rect 1660 693 1664 697
rect -68 662 2199 664
rect -4 661 2199 662
rect -4 658 1624 661
rect -68 657 1624 658
rect 1628 657 2199 661
rect -68 656 2199 657
rect 2479 662 2736 664
rect 2479 658 2672 662
rect 2479 656 2736 658
rect 1668 647 1672 651
rect -140 642 2199 644
rect -76 638 2199 642
rect -140 636 2199 638
rect 2479 642 2664 644
rect 2479 638 2600 642
rect 2479 636 2664 638
rect 856 596 875 600
rect 177 592 200 596
rect 361 592 384 596
rect 545 592 552 596
rect 705 592 712 596
rect 856 593 860 596
rect 1808 595 1812 599
rect 1801 591 1812 595
rect 2032 592 2067 596
rect 2032 588 2036 592
rect 1660 583 1664 587
rect -68 552 2199 554
rect -4 551 2199 552
rect -4 548 1624 551
rect -68 547 1624 548
rect 1628 547 2199 551
rect -68 546 2199 547
rect 2479 552 2736 554
rect 2479 548 2672 552
rect 2479 546 2736 548
rect 1668 537 1672 541
rect -140 532 2199 534
rect -76 528 2199 532
rect -140 526 2199 528
rect 2479 532 2664 534
rect 2479 528 2600 532
rect 2479 526 2664 528
rect 856 486 875 490
rect 177 482 208 486
rect 545 482 560 486
rect 705 482 720 486
rect 856 483 860 486
rect 1808 485 1812 489
rect 1801 481 1812 485
rect 2032 482 2067 486
rect 2032 478 2036 482
rect 1660 473 1664 477
rect -68 442 2199 444
rect -4 441 2199 442
rect -4 438 1624 441
rect -68 437 1624 438
rect 1628 437 2199 441
rect -68 436 2199 437
rect 2479 442 2736 444
rect 2479 438 2672 442
rect 2479 436 2736 438
rect 1668 427 1672 431
rect -140 422 2199 424
rect -76 418 2199 422
rect -140 416 2199 418
rect 2479 422 2664 424
rect 2479 418 2600 422
rect 2479 416 2664 418
rect 856 376 875 380
rect 177 372 216 376
rect 545 372 568 376
rect 705 372 728 376
rect 856 373 860 376
rect 1808 375 1812 379
rect 1801 371 1812 375
rect 2032 372 2067 376
rect 2032 368 2036 372
rect 1660 363 1664 367
rect -68 333 581 334
rect 758 333 2199 334
rect -68 332 2199 333
rect -4 331 2199 332
rect -4 328 1624 331
rect -68 327 1624 328
rect 1628 327 2199 331
rect -68 326 2199 327
rect 2479 332 2736 334
rect 2479 328 2672 332
rect 2479 326 2736 328
rect 573 325 925 326
rect 1668 317 1672 321
rect -140 312 2199 314
rect -76 308 2199 312
rect -140 306 2199 308
rect 2479 312 2664 314
rect 2479 308 2600 312
rect 2479 306 2664 308
rect 856 266 875 270
rect 177 262 224 266
rect 361 262 392 266
rect 705 262 736 266
rect 856 263 860 266
rect 1808 265 1812 269
rect 1801 261 1812 265
rect 2032 262 2067 266
rect 2032 258 2036 262
rect 1660 253 1664 257
rect -68 222 2199 224
rect -4 221 2199 222
rect -4 218 1624 221
rect -68 217 1624 218
rect 1628 217 2199 221
rect -68 216 2199 217
rect 2479 222 2736 224
rect 2479 218 2672 222
rect 2479 216 2736 218
rect 1668 207 1672 211
rect 2559 204 2563 206
rect -140 202 2199 204
rect -76 198 2199 202
rect 2479 202 2664 204
rect 2479 198 2600 202
rect -140 196 2197 198
rect 2479 196 2480 198
rect 2518 196 2522 198
rect 2545 196 2549 198
rect 2560 196 2664 198
rect 856 156 875 160
rect 361 152 400 156
rect 704 152 744 156
rect 856 153 860 156
rect 1808 155 1812 159
rect 1801 151 1812 155
rect 2032 152 2067 156
rect 2032 148 2036 152
rect -68 112 2199 114
rect -4 111 2199 112
rect -4 108 1624 111
rect -68 107 1624 108
rect 1628 107 1672 111
rect 1676 107 2199 111
rect -68 106 2199 107
rect 2479 112 2736 114
rect 2479 108 2672 112
rect 2479 106 2736 108
rect -140 92 2199 94
rect -76 91 2199 92
rect -76 88 1624 91
rect -140 87 1624 88
rect 1628 87 2199 91
rect -140 86 2199 87
rect 2479 92 2664 94
rect 2479 88 2600 92
rect 2479 86 2664 88
rect 856 46 875 50
rect 361 42 408 46
rect 704 42 752 46
rect 856 43 860 46
rect 1808 45 1812 49
rect 1801 41 1812 45
rect 2032 42 2067 46
rect 2032 38 2036 42
rect 1660 33 1664 37
rect -68 2 2199 4
rect -4 1 2199 2
rect -4 -2 1672 1
rect -68 -3 1672 -2
rect 1676 -3 2199 1
rect -68 -4 2199 -3
rect 2479 2 2736 4
rect 2479 -2 2672 2
rect 2479 -4 2736 -2
rect 2468 -252 2664 -248
rect 2468 -259 2600 -252
rect 2468 -263 2664 -259
rect -140 -276 949 -274
rect -76 -280 949 -276
rect -140 -282 949 -280
rect 2442 -277 2736 -273
rect 2442 -284 2672 -277
rect 2442 -289 2736 -284
rect -68 -366 948 -364
rect -4 -370 948 -366
rect -68 -372 948 -370
rect -140 -388 949 -386
rect -76 -392 949 -388
rect -140 -394 949 -392
rect -68 -478 952 -476
rect -4 -482 952 -478
rect -68 -484 950 -482
<< m2contact >>
rect -140 1298 -76 1302
rect 2600 1298 2664 1302
rect -68 1208 -4 1212
rect 2672 1208 2736 1212
rect 816 1198 820 1202
rect 856 1198 860 1202
rect 872 1198 876 1202
rect 888 1198 892 1202
rect -140 1188 -76 1192
rect 2600 1188 2664 1192
rect -68 1098 -4 1102
rect 2672 1098 2736 1102
rect 816 1088 820 1092
rect 872 1088 876 1092
rect -140 1078 -76 1082
rect 2600 1078 2664 1082
rect -68 988 -4 992
rect 2672 988 2736 992
rect -140 968 -76 972
rect 2600 968 2664 972
rect -68 878 -4 882
rect 2672 878 2736 882
rect -140 858 -76 862
rect 2600 858 2664 862
rect 184 812 188 816
rect 368 812 372 816
rect -68 768 -4 772
rect 1624 767 1628 771
rect 2672 768 2736 772
rect 1664 757 1668 761
rect 1672 757 1676 761
rect -140 748 -76 752
rect 2600 748 2664 752
rect 192 702 196 706
rect 376 702 380 706
rect 1656 693 1660 697
rect 1664 693 1668 697
rect -68 658 -4 662
rect 1624 657 1628 661
rect 2672 658 2736 662
rect 1664 647 1668 651
rect 1672 647 1676 651
rect -140 638 -76 642
rect 2600 638 2664 642
rect 200 592 204 596
rect 384 592 388 596
rect 552 592 556 596
rect 712 592 716 596
rect 1656 583 1660 587
rect 1664 583 1668 587
rect -68 548 -4 552
rect 1624 547 1628 551
rect 2672 548 2736 552
rect 1664 537 1668 541
rect 1672 537 1676 541
rect -140 528 -76 532
rect 2600 528 2664 532
rect 208 482 212 486
rect 560 482 564 486
rect 720 482 724 486
rect 1656 473 1660 477
rect 1664 473 1668 477
rect -68 438 -4 442
rect 1624 437 1628 441
rect 2672 438 2736 442
rect 1664 427 1668 431
rect 1672 427 1676 431
rect -140 418 -76 422
rect 2600 418 2664 422
rect 216 372 220 376
rect 568 372 572 376
rect 728 372 732 376
rect 1656 363 1660 367
rect 1664 363 1668 367
rect -68 328 -4 332
rect 1624 327 1628 331
rect 2672 328 2736 332
rect 1664 317 1668 321
rect 1672 317 1676 321
rect -140 308 -76 312
rect 2600 308 2664 312
rect 224 262 228 266
rect 392 262 396 266
rect 736 262 740 266
rect 1656 253 1660 257
rect 1664 253 1668 257
rect -68 218 -4 222
rect 1624 217 1628 221
rect 2672 218 2736 222
rect 1664 207 1668 211
rect 1672 207 1676 211
rect -140 198 -76 202
rect 2600 198 2664 202
rect 400 152 404 156
rect 744 152 748 156
rect -68 108 -4 112
rect 1624 107 1628 111
rect 1672 107 1676 111
rect 2672 108 2736 112
rect -140 88 -76 92
rect 1624 87 1628 91
rect 2600 88 2664 92
rect 408 42 412 46
rect 752 42 756 46
rect 1656 33 1660 37
rect 1664 33 1668 37
rect -68 -2 -4 2
rect 1672 -3 1676 1
rect 2672 -2 2736 2
rect 2600 -259 2664 -252
rect -140 -280 -76 -276
rect 2672 -284 2736 -277
rect -68 -370 -4 -366
rect -140 -392 -76 -388
rect -68 -482 -4 -478
<< metal2 >>
rect -140 1302 -76 1342
rect -140 1192 -76 1298
rect -140 1082 -76 1188
rect -140 972 -76 1078
rect -140 862 -76 968
rect -140 752 -76 858
rect -140 642 -76 748
rect -140 532 -76 638
rect -140 422 -76 528
rect -140 312 -76 418
rect -140 202 -76 308
rect -140 92 -76 198
rect -140 -276 -76 88
rect -140 -388 -76 -280
rect -140 -399 -76 -392
rect -68 1212 -4 1342
rect -68 1102 -4 1208
rect -68 992 -4 1098
rect -68 882 -4 988
rect 0 918 4 1312
rect 8 1203 12 1312
rect 16 1243 20 1312
rect 15 1242 21 1243
rect 15 1238 16 1242
rect 20 1238 21 1242
rect 15 1237 21 1238
rect 24 1223 28 1312
rect 23 1222 29 1223
rect 23 1218 24 1222
rect 28 1218 29 1222
rect 23 1217 29 1218
rect 7 1202 13 1203
rect 7 1198 8 1202
rect 12 1198 13 1202
rect 7 1197 13 1198
rect 56 918 60 1312
rect 135 1242 141 1243
rect 135 1238 136 1242
rect 140 1238 141 1242
rect 135 1237 141 1238
rect 136 963 140 1237
rect 135 962 141 963
rect 135 958 136 962
rect 140 958 141 962
rect 135 957 141 958
rect 87 952 93 953
rect 87 948 88 952
rect 92 948 93 952
rect 87 947 93 948
rect 88 939 92 947
rect 136 939 140 957
rect -68 772 -4 878
rect 63 852 69 853
rect 63 848 64 852
rect 68 848 69 852
rect 63 847 69 848
rect 39 832 45 833
rect 39 828 40 832
rect 44 828 45 832
rect 39 827 45 828
rect 0 813 4 819
rect -1 812 5 813
rect -1 808 0 812
rect 4 808 5 812
rect -1 807 5 808
rect 32 803 36 818
rect 40 808 44 827
rect 64 813 68 847
rect 184 816 188 1312
rect 31 802 37 803
rect 31 798 32 802
rect 36 798 37 802
rect 31 797 37 798
rect -68 662 -4 768
rect 63 742 69 743
rect 63 738 64 742
rect 68 738 69 742
rect 63 737 69 738
rect 39 722 45 723
rect 39 718 40 722
rect 44 718 45 722
rect 39 717 45 718
rect 0 703 4 709
rect -1 702 5 703
rect -1 698 0 702
rect 4 698 5 702
rect -1 697 5 698
rect 32 693 36 708
rect 40 698 44 717
rect 64 703 68 737
rect 192 706 196 1312
rect 31 692 37 693
rect 31 688 32 692
rect 36 688 37 692
rect 31 687 37 688
rect -68 552 -4 658
rect 63 632 69 633
rect 63 628 64 632
rect 68 628 69 632
rect 63 627 69 628
rect 39 612 45 613
rect 39 608 40 612
rect 44 608 45 612
rect 39 607 45 608
rect 0 593 4 599
rect -1 592 5 593
rect -1 588 0 592
rect 4 588 5 592
rect -1 587 5 588
rect 32 583 36 598
rect 40 588 44 607
rect 64 593 68 627
rect 200 596 204 1312
rect 31 582 37 583
rect 31 578 32 582
rect 36 578 37 582
rect 31 577 37 578
rect -68 442 -4 548
rect 63 522 69 523
rect 63 518 64 522
rect 68 518 69 522
rect 63 517 69 518
rect 39 502 45 503
rect 39 498 40 502
rect 44 498 45 502
rect 39 497 45 498
rect 0 483 4 489
rect -1 482 5 483
rect -1 478 0 482
rect 4 478 5 482
rect -1 477 5 478
rect 32 473 36 488
rect 40 478 44 497
rect 64 483 68 517
rect 208 486 212 1312
rect 31 472 37 473
rect 31 468 32 472
rect 36 468 37 472
rect 31 467 37 468
rect -68 332 -4 438
rect 63 412 69 413
rect 63 408 64 412
rect 68 408 69 412
rect 63 407 69 408
rect 39 392 45 393
rect 39 388 40 392
rect 44 388 45 392
rect 39 387 45 388
rect 0 373 4 379
rect -1 372 5 373
rect -1 368 0 372
rect 4 368 5 372
rect -1 367 5 368
rect 32 363 36 378
rect 40 368 44 387
rect 64 373 68 407
rect 216 376 220 1312
rect 31 362 37 363
rect 31 358 32 362
rect 36 358 37 362
rect 31 357 37 358
rect -68 222 -4 328
rect 63 302 69 303
rect 63 298 64 302
rect 68 298 69 302
rect 63 297 69 298
rect 39 282 45 283
rect 39 278 40 282
rect 44 278 45 282
rect 39 277 45 278
rect 0 263 4 269
rect -1 262 5 263
rect -1 258 0 262
rect 4 258 5 262
rect -1 257 5 258
rect 32 253 36 268
rect 40 258 44 277
rect 64 263 68 297
rect 224 266 228 1312
rect 240 918 244 1312
rect 391 1282 397 1283
rect 391 1278 392 1282
rect 396 1278 397 1282
rect 391 1277 397 1278
rect 392 1133 396 1277
rect 407 1182 413 1183
rect 407 1178 408 1182
rect 412 1178 413 1182
rect 407 1177 413 1178
rect 399 1172 405 1173
rect 399 1168 400 1172
rect 404 1168 405 1172
rect 399 1167 405 1168
rect 400 1163 404 1167
rect 399 1162 405 1163
rect 399 1158 400 1162
rect 404 1158 405 1162
rect 399 1157 405 1158
rect 391 1132 397 1133
rect 391 1128 392 1132
rect 396 1128 397 1132
rect 391 1127 397 1128
rect 383 1072 389 1073
rect 383 1068 384 1072
rect 388 1068 389 1072
rect 383 1067 389 1068
rect 375 1052 381 1053
rect 375 1048 376 1052
rect 380 1048 381 1052
rect 375 1047 381 1048
rect 367 1022 373 1023
rect 367 1018 368 1022
rect 372 1018 373 1022
rect 367 1017 373 1018
rect 319 962 325 963
rect 319 958 320 962
rect 324 958 325 962
rect 319 957 325 958
rect 271 952 277 953
rect 271 948 272 952
rect 276 948 277 952
rect 271 947 277 948
rect 272 939 276 947
rect 320 939 324 957
rect 247 852 253 853
rect 247 848 248 852
rect 252 848 253 852
rect 247 847 253 848
rect 248 813 252 847
rect 368 816 372 1017
rect 247 742 253 743
rect 247 738 248 742
rect 252 738 253 742
rect 247 737 253 738
rect 248 703 252 737
rect 376 706 380 1047
rect 247 632 253 633
rect 247 628 248 632
rect 252 628 253 632
rect 247 627 253 628
rect 248 593 252 627
rect 384 596 388 1067
rect 247 522 253 523
rect 247 518 248 522
rect 252 518 253 522
rect 247 517 253 518
rect 248 483 252 517
rect 247 412 253 413
rect 247 408 248 412
rect 252 408 253 412
rect 247 407 253 408
rect 248 373 252 407
rect 247 302 253 303
rect 247 298 248 302
rect 252 298 253 302
rect 247 297 253 298
rect 248 263 252 297
rect 392 266 396 1127
rect 31 252 37 253
rect 31 248 32 252
rect 36 248 37 252
rect 31 247 37 248
rect -68 112 -4 218
rect 63 192 69 193
rect 63 188 64 192
rect 68 188 69 192
rect 63 187 69 188
rect 247 192 253 193
rect 247 188 248 192
rect 252 188 253 192
rect 247 187 253 188
rect 39 172 45 173
rect 39 168 40 172
rect 44 168 45 172
rect 39 167 45 168
rect 0 153 4 159
rect -1 152 5 153
rect -1 148 0 152
rect 4 148 5 152
rect -1 147 5 148
rect 32 143 36 158
rect 40 148 44 167
rect 64 153 68 187
rect 248 153 252 187
rect 400 156 404 1157
rect 408 1063 412 1177
rect 407 1062 413 1063
rect 407 1058 408 1062
rect 412 1058 413 1062
rect 407 1057 413 1058
rect 31 142 37 143
rect 31 138 32 142
rect 36 138 37 142
rect 31 137 37 138
rect -68 2 -4 108
rect 63 82 69 83
rect 63 78 64 82
rect 68 78 69 82
rect 63 77 69 78
rect 247 82 253 83
rect 247 78 248 82
rect 252 78 253 82
rect 247 77 253 78
rect 39 62 45 63
rect 39 58 40 62
rect 44 58 45 62
rect 39 57 45 58
rect 0 43 4 49
rect -1 42 5 43
rect -1 38 0 42
rect 4 38 5 42
rect -1 37 5 38
rect 32 33 36 48
rect 40 38 44 57
rect 64 43 68 77
rect 248 43 252 77
rect 408 46 412 1057
rect 424 918 428 1312
rect 551 1262 557 1263
rect 551 1258 552 1262
rect 556 1258 557 1262
rect 551 1257 557 1258
rect 503 962 509 963
rect 503 958 504 962
rect 508 958 509 962
rect 503 957 509 958
rect 455 952 461 953
rect 455 948 456 952
rect 460 948 461 952
rect 455 947 461 948
rect 456 939 460 947
rect 504 939 508 957
rect 431 852 437 853
rect 431 848 432 852
rect 436 848 437 852
rect 431 847 437 848
rect 432 813 436 847
rect 431 742 437 743
rect 431 738 432 742
rect 436 738 437 742
rect 431 737 437 738
rect 432 703 436 737
rect 431 632 437 633
rect 431 628 432 632
rect 436 628 437 632
rect 431 627 437 628
rect 432 593 436 627
rect 552 596 556 1257
rect 559 1152 565 1153
rect 559 1148 560 1152
rect 564 1148 565 1152
rect 559 1147 565 1148
rect 431 522 437 523
rect 431 518 432 522
rect 436 518 437 522
rect 431 517 437 518
rect 432 483 436 517
rect 560 486 564 1147
rect 567 1042 573 1043
rect 567 1038 568 1042
rect 572 1038 573 1042
rect 567 1037 573 1038
rect 431 412 437 413
rect 431 408 432 412
rect 436 408 437 412
rect 431 407 437 408
rect 432 373 436 407
rect 568 376 572 1037
rect 584 918 588 1312
rect 615 1222 621 1223
rect 615 1218 616 1222
rect 620 1218 621 1222
rect 615 1217 621 1218
rect 616 953 620 1217
rect 663 962 669 963
rect 663 958 664 962
rect 668 958 669 962
rect 663 957 669 958
rect 615 952 621 953
rect 615 948 616 952
rect 620 948 621 952
rect 615 947 621 948
rect 616 939 620 947
rect 664 939 668 957
rect 696 943 700 1312
rect 695 942 701 943
rect 695 938 696 942
rect 700 938 701 942
rect 695 937 701 938
rect 591 852 597 853
rect 591 848 592 852
rect 596 848 597 852
rect 591 847 597 848
rect 592 813 596 847
rect 703 832 709 833
rect 591 742 597 743
rect 591 738 592 742
rect 596 738 597 742
rect 591 737 597 738
rect 592 703 596 737
rect 591 632 597 633
rect 591 628 592 632
rect 596 628 597 632
rect 591 627 597 628
rect 592 593 596 627
rect 591 522 597 523
rect 591 518 592 522
rect 596 518 597 522
rect 591 517 597 518
rect 592 483 596 517
rect 591 412 597 413
rect 591 408 592 412
rect 596 408 597 412
rect 591 407 597 408
rect 592 373 596 407
rect 431 302 437 303
rect 431 298 432 302
rect 436 298 437 302
rect 431 297 437 298
rect 591 302 597 303
rect 591 298 592 302
rect 596 298 597 302
rect 591 297 597 298
rect 432 263 436 297
rect 592 263 596 297
rect 431 192 437 193
rect 431 188 432 192
rect 436 188 437 192
rect 431 187 437 188
rect 591 192 597 193
rect 591 188 592 192
rect 596 188 597 192
rect 591 187 597 188
rect 432 153 436 187
rect 592 153 596 187
rect 431 82 437 83
rect 431 78 432 82
rect 436 78 437 82
rect 431 77 437 78
rect 591 82 597 83
rect 591 78 592 82
rect 596 78 597 82
rect 591 77 597 78
rect 432 43 436 77
rect 31 32 37 33
rect 31 28 32 32
rect 36 28 37 32
rect 31 27 37 28
rect -68 -366 -4 -2
rect 544 -152 548 46
rect 592 43 596 77
rect 617 -170 621 718
rect 696 -161 700 828
rect 703 828 704 832
rect 708 828 709 832
rect 703 827 709 828
rect 704 812 708 827
rect 703 722 709 723
rect 703 718 704 722
rect 708 718 709 722
rect 703 717 709 718
rect 704 702 708 717
rect 703 612 709 613
rect 703 608 704 612
rect 708 608 709 612
rect 703 607 709 608
rect 704 592 708 607
rect 712 596 716 1312
rect 703 502 709 503
rect 703 498 704 502
rect 708 498 709 502
rect 703 497 709 498
rect 704 482 708 497
rect 720 486 724 1312
rect 703 392 709 393
rect 703 388 704 392
rect 708 388 709 392
rect 703 387 709 388
rect 704 372 708 387
rect 728 376 732 1312
rect 703 282 709 283
rect 703 278 704 282
rect 708 278 709 282
rect 703 277 709 278
rect 704 262 708 277
rect 736 266 740 1312
rect 703 172 709 173
rect 703 168 704 172
rect 708 168 709 172
rect 703 167 709 168
rect 704 152 708 167
rect 744 156 748 1312
rect 703 62 709 63
rect 703 58 704 62
rect 708 58 709 62
rect 703 57 709 58
rect 704 42 708 57
rect 752 46 756 1312
rect 767 1262 773 1263
rect 767 1258 768 1262
rect 772 1258 773 1262
rect 767 1257 773 1258
rect 768 1254 772 1257
rect 767 1152 773 1153
rect 767 1148 768 1152
rect 772 1148 773 1152
rect 767 1147 773 1148
rect 768 1144 772 1147
rect 767 1042 773 1043
rect 767 1038 768 1042
rect 772 1038 773 1042
rect 792 1041 796 1312
rect 799 1282 805 1283
rect 799 1278 800 1282
rect 804 1278 805 1282
rect 799 1277 805 1278
rect 800 1264 804 1277
rect 856 1202 860 1251
rect 888 1202 892 1251
rect 960 1248 964 1312
rect 1496 1293 1500 1312
rect 799 1172 805 1173
rect 799 1168 800 1172
rect 804 1168 805 1172
rect 799 1167 805 1168
rect 800 1154 804 1167
rect 816 1139 820 1198
rect 872 1092 876 1198
rect 799 1062 805 1063
rect 799 1058 800 1062
rect 804 1058 805 1062
rect 799 1057 805 1058
rect 800 1044 804 1057
rect 767 1037 773 1038
rect 768 1034 772 1037
rect 816 1029 820 1088
rect 815 962 821 963
rect 815 958 816 962
rect 820 958 821 962
rect 815 957 821 958
rect 767 952 773 953
rect 767 948 768 952
rect 772 948 773 952
rect 767 947 773 948
rect 768 939 772 947
rect 816 939 820 957
rect 871 942 877 943
rect 871 938 872 942
rect 876 938 877 942
rect 871 937 877 938
rect 872 919 876 937
rect 767 852 773 853
rect 767 848 768 852
rect 772 848 773 852
rect 767 847 773 848
rect 768 813 772 847
rect 911 822 917 823
rect 911 818 912 822
rect 916 818 917 822
rect 911 817 917 818
rect 904 813 908 817
rect 903 812 909 813
rect 903 808 904 812
rect 908 808 909 812
rect 912 809 916 817
rect 903 807 909 808
rect 767 742 773 743
rect 767 738 768 742
rect 772 738 773 742
rect 767 737 773 738
rect 768 703 772 737
rect 911 712 917 713
rect 911 708 912 712
rect 916 708 917 712
rect 911 707 917 708
rect 904 703 908 707
rect 903 702 909 703
rect 903 698 904 702
rect 908 698 909 702
rect 912 699 916 707
rect 903 697 909 698
rect 767 632 773 633
rect 767 628 768 632
rect 772 628 773 632
rect 767 627 773 628
rect 768 593 772 627
rect 911 602 917 603
rect 911 598 912 602
rect 916 598 917 602
rect 911 597 917 598
rect 904 593 908 597
rect 903 592 909 593
rect 903 588 904 592
rect 908 588 909 592
rect 912 589 916 597
rect 903 587 909 588
rect 767 522 773 523
rect 767 518 768 522
rect 772 518 773 522
rect 767 517 773 518
rect 768 483 772 517
rect 911 492 917 493
rect 911 488 912 492
rect 916 488 917 492
rect 911 487 917 488
rect 904 483 908 487
rect 903 482 909 483
rect 903 478 904 482
rect 908 478 909 482
rect 912 479 916 487
rect 903 477 909 478
rect 767 412 773 413
rect 767 408 768 412
rect 772 408 773 412
rect 767 407 773 408
rect 768 373 772 407
rect 911 382 917 383
rect 911 378 912 382
rect 916 378 917 382
rect 911 377 917 378
rect 904 373 908 377
rect 903 372 909 373
rect 903 368 904 372
rect 908 368 909 372
rect 912 369 916 377
rect 903 367 909 368
rect 767 302 773 303
rect 767 298 768 302
rect 772 298 773 302
rect 767 297 773 298
rect 768 263 772 297
rect 911 272 917 273
rect 911 268 912 272
rect 916 268 917 272
rect 911 267 917 268
rect 904 263 908 267
rect 903 262 909 263
rect 903 258 904 262
rect 908 258 909 262
rect 912 259 916 267
rect 903 257 909 258
rect 767 192 773 193
rect 767 188 768 192
rect 772 188 773 192
rect 767 187 773 188
rect 768 153 772 187
rect 911 162 917 163
rect 911 158 912 162
rect 916 158 917 162
rect 911 157 917 158
rect 904 153 908 157
rect 903 152 909 153
rect 903 148 904 152
rect 908 148 909 152
rect 912 149 916 157
rect 903 147 909 148
rect 767 82 773 83
rect 767 78 768 82
rect 772 78 773 82
rect 767 77 773 78
rect 768 43 772 77
rect 911 52 917 53
rect 911 48 912 52
rect 916 48 917 52
rect 911 47 917 48
rect 904 43 908 47
rect 903 42 909 43
rect 903 38 904 42
rect 908 38 909 42
rect 912 39 916 47
rect 903 37 909 38
rect 998 -187 1002 -66
rect 1078 -184 1082 -57
rect 1158 -185 1162 -48
rect 1190 -184 1194 -75
rect 1238 -184 1242 -39
rect 1318 -184 1322 -30
rect 1398 -185 1402 -21
rect 1478 -185 1482 -12
rect 1496 -183 1500 1289
rect 1584 1284 1588 1312
rect 1551 962 1557 963
rect 1551 958 1552 962
rect 1556 958 1557 962
rect 1551 957 1557 958
rect 1503 952 1509 953
rect 1503 948 1504 952
rect 1508 948 1509 952
rect 1503 947 1509 948
rect 1504 939 1508 947
rect 1552 939 1556 957
rect 1504 783 1508 816
rect 1503 782 1509 783
rect 1503 778 1504 782
rect 1508 778 1509 782
rect 1503 777 1509 778
rect 1504 673 1508 706
rect 1503 672 1509 673
rect 1503 668 1504 672
rect 1508 668 1509 672
rect 1503 667 1509 668
rect 1504 563 1508 596
rect 1503 562 1509 563
rect 1503 558 1504 562
rect 1508 558 1509 562
rect 1503 557 1509 558
rect 1504 453 1508 486
rect 1503 452 1509 453
rect 1503 448 1504 452
rect 1508 448 1509 452
rect 1503 447 1509 448
rect 1504 343 1508 376
rect 1503 342 1509 343
rect 1503 338 1504 342
rect 1508 338 1509 342
rect 1503 337 1509 338
rect 1504 233 1508 266
rect 1503 232 1509 233
rect 1503 228 1504 232
rect 1508 228 1509 232
rect 1503 227 1509 228
rect 1504 123 1508 156
rect 1503 122 1509 123
rect 1503 118 1504 122
rect 1508 118 1509 122
rect 1503 117 1509 118
rect 1504 13 1508 46
rect 1503 12 1509 13
rect 1503 8 1504 12
rect 1508 8 1509 12
rect 1503 7 1509 8
rect 1584 2 1588 1280
rect 1600 918 1604 1312
rect 1632 918 1636 1312
rect 1759 962 1765 963
rect 1759 958 1760 962
rect 1764 958 1765 962
rect 1759 957 1765 958
rect 1711 952 1717 953
rect 1711 948 1712 952
rect 1716 948 1717 952
rect 1711 947 1717 948
rect 1712 939 1716 947
rect 1760 939 1764 957
rect 1808 918 1812 1312
rect 1911 962 1917 963
rect 1911 958 1912 962
rect 1916 958 1917 962
rect 1911 957 1917 958
rect 1863 952 1869 953
rect 1863 948 1864 952
rect 1868 948 1869 952
rect 1863 947 1869 948
rect 1864 939 1868 947
rect 1912 939 1916 957
rect 1960 918 1964 1312
rect 1992 918 1996 1312
rect 2048 918 2052 1312
rect 2079 1202 2085 1203
rect 2079 1198 2080 1202
rect 2084 1198 2085 1202
rect 2079 1197 2085 1198
rect 2080 918 2084 1197
rect 2143 962 2149 963
rect 2143 958 2144 962
rect 2148 958 2149 962
rect 2143 957 2149 958
rect 2095 952 2101 953
rect 2095 948 2096 952
rect 2100 948 2101 952
rect 2095 947 2101 948
rect 2096 939 2100 947
rect 2144 939 2148 957
rect 2186 852 2190 853
rect 1847 851 1853 852
rect 1847 847 1848 851
rect 1852 847 1853 851
rect 1847 846 1853 847
rect 1591 842 1597 843
rect 1591 838 1592 842
rect 1596 838 1597 842
rect 1591 837 1597 838
rect 1615 842 1621 843
rect 1615 838 1616 842
rect 1620 838 1621 842
rect 1615 837 1621 838
rect 1695 842 1701 843
rect 1695 838 1696 842
rect 1700 838 1701 842
rect 1695 837 1701 838
rect 1592 812 1596 837
rect 1616 804 1620 837
rect 1655 832 1661 833
rect 1655 828 1656 832
rect 1660 828 1661 832
rect 1655 827 1661 828
rect 1671 832 1677 833
rect 1671 828 1672 832
rect 1676 828 1677 832
rect 1671 827 1677 828
rect 1656 819 1660 827
rect 1624 771 1628 807
rect 1672 761 1676 827
rect 1696 807 1700 837
rect 1712 793 1716 816
rect 1840 803 1844 818
rect 1848 808 1852 846
rect 2015 832 2021 833
rect 2015 828 2016 832
rect 2020 828 2021 832
rect 2015 827 2021 828
rect 1839 802 1845 803
rect 1839 798 1840 802
rect 1844 798 1845 802
rect 1839 797 1845 798
rect 1711 792 1717 793
rect 1711 788 1712 792
rect 1716 788 1717 792
rect 1711 787 1717 788
rect 1864 783 1868 816
rect 1952 813 1956 815
rect 1976 813 1980 821
rect 2016 818 2020 827
rect 1951 812 1957 813
rect 1975 812 1981 813
rect 1951 808 1952 812
rect 1956 808 1957 812
rect 1951 807 1957 808
rect 1968 783 1972 812
rect 1975 808 1976 812
rect 1980 808 1981 812
rect 1975 807 1981 808
rect 1863 782 1869 783
rect 1863 778 1864 782
rect 1868 778 1869 782
rect 1863 777 1869 778
rect 1967 782 1973 783
rect 1967 778 1968 782
rect 1972 778 1973 782
rect 1967 777 1973 778
rect 1591 732 1597 733
rect 1591 728 1592 732
rect 1596 728 1597 732
rect 1591 727 1597 728
rect 1615 732 1621 733
rect 1615 728 1616 732
rect 1620 728 1621 732
rect 1615 727 1621 728
rect 1592 702 1596 727
rect 1616 694 1620 727
rect 1655 722 1661 723
rect 1655 718 1656 722
rect 1660 718 1661 722
rect 1655 717 1661 718
rect 1656 709 1660 717
rect 1664 697 1668 757
rect 2168 752 2172 838
rect 2176 830 2180 838
rect 2186 817 2190 848
rect 2176 803 2180 812
rect 2175 802 2181 803
rect 2175 798 2176 802
rect 2180 798 2181 802
rect 2175 797 2181 798
rect 2176 762 2180 778
rect 2176 757 2180 758
rect 1671 722 1677 723
rect 1671 718 1672 722
rect 1676 718 1677 722
rect 1671 717 1677 718
rect 1624 661 1628 697
rect 1591 622 1597 623
rect 1591 618 1592 622
rect 1596 618 1597 622
rect 1591 617 1597 618
rect 1615 622 1621 623
rect 1615 618 1616 622
rect 1620 618 1621 622
rect 1615 617 1621 618
rect 1592 592 1596 617
rect 1616 584 1620 617
rect 1656 613 1660 693
rect 1672 651 1676 717
rect 1655 612 1661 613
rect 1655 608 1656 612
rect 1660 608 1661 612
rect 1655 607 1661 608
rect 1656 599 1660 607
rect 1664 587 1668 647
rect 1671 612 1677 613
rect 1671 608 1672 612
rect 1676 608 1677 612
rect 1671 607 1677 608
rect 1624 551 1628 587
rect 1591 512 1597 513
rect 1591 508 1592 512
rect 1596 508 1597 512
rect 1591 507 1597 508
rect 1615 512 1621 513
rect 1615 508 1616 512
rect 1620 508 1621 512
rect 1615 507 1621 508
rect 1592 482 1596 507
rect 1616 474 1620 507
rect 1656 503 1660 583
rect 1672 541 1676 607
rect 1655 502 1661 503
rect 1655 498 1656 502
rect 1660 498 1661 502
rect 1655 497 1661 498
rect 1656 489 1660 497
rect 1664 477 1668 537
rect 1671 502 1677 503
rect 1671 498 1672 502
rect 1676 498 1677 502
rect 1671 497 1677 498
rect 1624 441 1628 477
rect 1591 402 1597 403
rect 1591 398 1592 402
rect 1596 398 1597 402
rect 1591 397 1597 398
rect 1615 402 1621 403
rect 1615 398 1616 402
rect 1620 398 1621 402
rect 1615 397 1621 398
rect 1592 372 1596 397
rect 1616 364 1620 397
rect 1656 393 1660 473
rect 1672 431 1676 497
rect 1655 392 1661 393
rect 1655 388 1656 392
rect 1660 388 1661 392
rect 1655 387 1661 388
rect 1656 379 1660 387
rect 1664 367 1668 427
rect 1671 392 1677 393
rect 1671 388 1672 392
rect 1676 388 1677 392
rect 1671 387 1677 388
rect 1624 331 1628 367
rect 1591 292 1597 293
rect 1591 288 1592 292
rect 1596 288 1597 292
rect 1591 287 1597 288
rect 1615 292 1621 293
rect 1615 288 1616 292
rect 1620 288 1621 292
rect 1615 287 1621 288
rect 1592 262 1596 287
rect 1616 254 1620 287
rect 1656 283 1660 363
rect 1672 321 1676 387
rect 1655 282 1661 283
rect 1655 278 1656 282
rect 1660 278 1661 282
rect 1655 277 1661 278
rect 1656 269 1660 277
rect 1664 257 1668 317
rect 1671 282 1677 283
rect 1671 278 1672 282
rect 1676 278 1677 282
rect 1671 277 1677 278
rect 1624 221 1628 257
rect 1591 182 1597 183
rect 1591 178 1592 182
rect 1596 178 1597 182
rect 1591 177 1597 178
rect 1615 182 1621 183
rect 1615 178 1616 182
rect 1620 178 1621 182
rect 1615 177 1621 178
rect 1592 152 1596 177
rect 1616 144 1620 177
rect 1656 173 1660 253
rect 1672 211 1676 277
rect 1655 172 1661 173
rect 1655 168 1656 172
rect 1660 168 1661 172
rect 1655 167 1661 168
rect 1656 159 1660 167
rect 1624 111 1628 147
rect 1591 72 1597 73
rect 1591 68 1592 72
rect 1596 68 1597 72
rect 1591 67 1597 68
rect 1615 72 1621 73
rect 1615 68 1616 72
rect 1620 68 1621 72
rect 1615 67 1621 68
rect 1592 42 1596 67
rect 1616 34 1620 67
rect 1624 34 1628 87
rect 1655 62 1661 63
rect 1655 58 1656 62
rect 1660 58 1661 62
rect 1655 57 1661 58
rect 1656 37 1660 57
rect 1664 37 1668 207
rect 1671 172 1677 173
rect 1671 168 1672 172
rect 1676 168 1677 172
rect 1671 167 1677 168
rect 1672 111 1676 167
rect 1671 62 1677 63
rect 1671 58 1672 62
rect 1676 58 1677 62
rect 1671 57 1677 58
rect 1672 1 1676 57
rect 1529 -185 1533 -2
rect 1688 -8 1692 748
rect 2186 742 2190 743
rect 1847 741 1853 742
rect 1847 737 1848 741
rect 1852 737 1853 741
rect 1847 736 1853 737
rect 1695 732 1701 733
rect 1695 728 1696 732
rect 1700 728 1701 732
rect 1695 727 1701 728
rect 1696 697 1700 727
rect 1712 683 1716 706
rect 1840 693 1844 708
rect 1848 698 1852 736
rect 2015 722 2021 723
rect 2015 718 2016 722
rect 2020 718 2021 722
rect 2015 717 2021 718
rect 1839 692 1845 693
rect 1839 688 1840 692
rect 1844 688 1845 692
rect 1839 687 1845 688
rect 1711 682 1717 683
rect 1711 678 1712 682
rect 1716 678 1717 682
rect 1711 677 1717 678
rect 1864 673 1868 706
rect 1952 703 1956 705
rect 1976 703 1980 711
rect 2016 708 2020 717
rect 1951 702 1957 703
rect 1975 702 1981 703
rect 1951 698 1952 702
rect 1956 698 1957 702
rect 1951 697 1957 698
rect 1968 673 1972 702
rect 1975 698 1976 702
rect 1980 698 1981 702
rect 1975 697 1981 698
rect 1863 672 1869 673
rect 1863 668 1864 672
rect 1868 668 1869 672
rect 1863 667 1869 668
rect 1967 672 1973 673
rect 1967 668 1968 672
rect 1972 668 1973 672
rect 1967 667 1973 668
rect 2168 642 2172 728
rect 2176 720 2180 728
rect 2186 707 2190 738
rect 2176 693 2180 702
rect 2175 692 2181 693
rect 2175 688 2176 692
rect 2180 688 2181 692
rect 2175 687 2181 688
rect 2176 652 2180 668
rect 2176 647 2180 648
rect 1695 622 1701 623
rect 1695 618 1696 622
rect 1700 618 1701 622
rect 1695 617 1701 618
rect 1696 587 1700 617
rect 1695 512 1701 513
rect 1695 508 1696 512
rect 1700 508 1701 512
rect 1695 507 1701 508
rect 1696 477 1700 507
rect 1695 402 1701 403
rect 1695 398 1696 402
rect 1700 398 1701 402
rect 1695 397 1701 398
rect 1696 367 1700 397
rect 1695 292 1701 293
rect 1695 288 1696 292
rect 1700 288 1701 292
rect 1695 287 1701 288
rect 1696 257 1700 287
rect 1695 182 1701 183
rect 1695 178 1696 182
rect 1700 178 1701 182
rect 1695 177 1701 178
rect 1696 147 1700 177
rect 1695 72 1701 73
rect 1695 68 1696 72
rect 1700 68 1701 72
rect 1695 67 1701 68
rect 1696 37 1700 67
rect 1704 -17 1708 638
rect 2186 632 2190 633
rect 1847 631 1853 632
rect 1847 627 1848 631
rect 1852 627 1853 631
rect 1847 626 1853 627
rect 1712 573 1716 596
rect 1840 583 1844 598
rect 1848 588 1852 626
rect 2015 612 2021 613
rect 2015 608 2016 612
rect 2020 608 2021 612
rect 2015 607 2021 608
rect 1839 582 1845 583
rect 1839 578 1840 582
rect 1844 578 1845 582
rect 1839 577 1845 578
rect 1711 572 1717 573
rect 1711 568 1712 572
rect 1716 568 1717 572
rect 1711 567 1717 568
rect 1864 563 1868 596
rect 1952 593 1956 595
rect 1976 593 1980 601
rect 2016 598 2020 607
rect 1951 592 1957 593
rect 1975 592 1981 593
rect 1951 588 1952 592
rect 1956 588 1957 592
rect 1951 587 1957 588
rect 1968 563 1972 592
rect 1975 588 1976 592
rect 1980 588 1981 592
rect 1975 587 1981 588
rect 1863 562 1869 563
rect 1863 558 1864 562
rect 1868 558 1869 562
rect 1863 557 1869 558
rect 1967 562 1973 563
rect 1967 558 1968 562
rect 1972 558 1973 562
rect 1967 557 1973 558
rect 2168 532 2172 618
rect 2176 610 2180 618
rect 2186 597 2190 628
rect 2176 583 2180 592
rect 2175 582 2181 583
rect 2175 578 2176 582
rect 2180 578 2181 582
rect 2175 577 2181 578
rect 2176 542 2180 558
rect 2176 537 2180 538
rect 1712 463 1716 486
rect 1711 462 1717 463
rect 1711 458 1712 462
rect 1716 458 1717 462
rect 1711 457 1717 458
rect 1712 353 1716 376
rect 1711 352 1717 353
rect 1711 348 1712 352
rect 1716 348 1717 352
rect 1711 347 1717 348
rect 1712 243 1716 266
rect 1711 242 1717 243
rect 1711 238 1712 242
rect 1716 238 1717 242
rect 1711 237 1717 238
rect 1712 133 1716 156
rect 1711 132 1717 133
rect 1711 128 1712 132
rect 1716 128 1717 132
rect 1711 127 1717 128
rect 1712 23 1716 46
rect 1711 22 1717 23
rect 1711 18 1712 22
rect 1716 18 1717 22
rect 1711 17 1717 18
rect 1792 -26 1796 528
rect 2186 522 2190 523
rect 1847 521 1853 522
rect 1847 517 1848 521
rect 1852 517 1853 521
rect 1847 516 1853 517
rect 1840 473 1844 488
rect 1848 478 1852 516
rect 2015 502 2021 503
rect 2015 498 2016 502
rect 2020 498 2021 502
rect 2015 497 2021 498
rect 1839 472 1845 473
rect 1839 468 1840 472
rect 1844 468 1845 472
rect 1839 467 1845 468
rect 1864 453 1868 486
rect 1952 483 1956 485
rect 1976 483 1980 491
rect 2016 488 2020 497
rect 1951 482 1957 483
rect 1975 482 1981 483
rect 1951 478 1952 482
rect 1956 478 1957 482
rect 1951 477 1957 478
rect 1968 453 1972 482
rect 1975 478 1976 482
rect 1980 478 1981 482
rect 1975 477 1981 478
rect 1863 452 1869 453
rect 1863 448 1864 452
rect 1868 448 1869 452
rect 1863 447 1869 448
rect 1967 452 1973 453
rect 1967 448 1968 452
rect 1972 448 1973 452
rect 1967 447 1973 448
rect 2168 422 2172 508
rect 2176 500 2180 508
rect 2186 487 2190 518
rect 2176 473 2180 482
rect 2175 472 2181 473
rect 2175 468 2176 472
rect 2180 468 2181 472
rect 2175 467 2181 468
rect 2176 432 2180 448
rect 2176 427 2180 428
rect 1847 411 1853 412
rect 1847 407 1848 411
rect 1852 407 1853 411
rect 1847 406 1853 407
rect 1840 363 1844 378
rect 1848 368 1852 406
rect 1839 362 1845 363
rect 1839 358 1840 362
rect 1844 358 1845 362
rect 1839 357 1845 358
rect 1847 301 1853 302
rect 1847 297 1848 301
rect 1852 297 1853 301
rect 1847 296 1853 297
rect 1840 253 1844 268
rect 1848 258 1852 296
rect 1839 252 1845 253
rect 1839 248 1840 252
rect 1844 248 1845 252
rect 1839 247 1845 248
rect 1847 191 1853 192
rect 1847 187 1848 191
rect 1852 187 1853 191
rect 1847 186 1853 187
rect 1840 143 1844 158
rect 1848 148 1852 186
rect 1839 142 1845 143
rect 1839 138 1840 142
rect 1844 138 1845 142
rect 1839 137 1845 138
rect 1847 81 1853 82
rect 1847 77 1848 81
rect 1852 77 1853 81
rect 1847 76 1853 77
rect 1840 33 1844 48
rect 1848 38 1852 76
rect 1839 32 1845 33
rect 1839 28 1840 32
rect 1844 28 1845 32
rect 1839 27 1845 28
rect 1856 -35 1860 418
rect 2015 392 2021 393
rect 2015 388 2016 392
rect 2020 388 2021 392
rect 2015 387 2021 388
rect 1864 343 1868 376
rect 1952 373 1956 375
rect 1976 373 1980 381
rect 2016 378 2020 387
rect 1951 372 1957 373
rect 1975 372 1981 373
rect 1951 368 1952 372
rect 1956 368 1957 372
rect 1951 367 1957 368
rect 1968 343 1972 372
rect 1975 368 1976 372
rect 1980 368 1981 372
rect 1975 367 1981 368
rect 1863 342 1869 343
rect 1863 338 1864 342
rect 1868 338 1869 342
rect 1863 337 1869 338
rect 1967 342 1973 343
rect 1967 338 1968 342
rect 1972 338 1973 342
rect 1967 337 1973 338
rect 2168 312 2172 398
rect 2176 390 2180 398
rect 2186 377 2190 413
rect 2176 363 2180 372
rect 2175 362 2181 363
rect 2175 358 2176 362
rect 2180 358 2181 362
rect 2175 357 2181 358
rect 2176 322 2180 338
rect 1864 233 1868 266
rect 1863 232 1869 233
rect 1863 228 1864 232
rect 1868 228 1869 232
rect 1863 227 1869 228
rect 1864 123 1868 156
rect 1863 122 1869 123
rect 1863 118 1864 122
rect 1868 118 1869 122
rect 1863 117 1869 118
rect 1864 13 1868 46
rect 1863 12 1869 13
rect 1863 8 1864 12
rect 1868 8 1869 12
rect 1863 7 1869 8
rect 1944 -44 1948 308
rect 2185 302 2189 303
rect 2015 282 2021 283
rect 2015 278 2016 282
rect 2020 278 2021 282
rect 2015 277 2021 278
rect 1952 263 1956 265
rect 1976 263 1980 271
rect 2016 268 2020 277
rect 1951 262 1957 263
rect 1975 262 1981 263
rect 1951 258 1952 262
rect 1956 258 1957 262
rect 1951 257 1957 258
rect 1968 233 1972 262
rect 1975 258 1976 262
rect 1980 258 1981 262
rect 1975 257 1981 258
rect 1967 232 1973 233
rect 1967 228 1968 232
rect 1972 228 1973 232
rect 1967 227 1973 228
rect 2168 202 2172 288
rect 2176 280 2180 288
rect 2185 267 2189 298
rect 2176 253 2180 262
rect 2175 252 2181 253
rect 2175 248 2176 252
rect 2180 248 2181 252
rect 2175 247 2181 248
rect 2176 212 2180 228
rect 1952 153 1956 155
rect 1976 153 1980 161
rect 1951 152 1957 153
rect 1975 152 1981 153
rect 1951 148 1952 152
rect 1956 148 1957 152
rect 1951 147 1957 148
rect 1968 123 1972 152
rect 1975 148 1976 152
rect 1980 148 1981 152
rect 1975 147 1981 148
rect 1967 122 1973 123
rect 1967 118 1968 122
rect 1972 118 1973 122
rect 1967 117 1973 118
rect 1952 43 1956 45
rect 1976 43 1980 51
rect 1951 42 1957 43
rect 1975 42 1981 43
rect 1951 38 1952 42
rect 1956 38 1957 42
rect 1951 37 1957 38
rect 1968 13 1972 42
rect 1975 38 1976 42
rect 1980 38 1981 42
rect 1975 37 1981 38
rect 1967 12 1973 13
rect 1967 8 1968 12
rect 1972 8 1973 12
rect 1967 7 1973 8
rect 1992 -53 1996 198
rect 2186 192 2190 193
rect 2015 172 2021 173
rect 2015 168 2016 172
rect 2020 168 2021 172
rect 2015 167 2021 168
rect 2016 158 2020 167
rect 2024 92 2028 93
rect 2168 92 2172 178
rect 2176 172 2180 178
rect 2186 159 2190 188
rect 2176 143 2180 152
rect 2175 142 2181 143
rect 2175 138 2176 142
rect 2180 138 2181 142
rect 2175 137 2181 138
rect 2176 102 2180 118
rect 2015 62 2021 63
rect 2015 58 2016 62
rect 2020 58 2021 62
rect 2015 57 2021 58
rect 2016 48 2020 57
rect 2024 -62 2028 88
rect 2186 82 2190 83
rect 2168 -71 2172 68
rect 2176 60 2180 68
rect 2186 47 2190 78
rect 2176 33 2180 42
rect 2175 32 2181 33
rect 2175 28 2176 32
rect 2180 28 2181 32
rect 2175 27 2181 28
rect 2176 -9 2180 8
rect 1544 -187 1548 -84
rect 1566 -186 1570 -93
rect 1588 -185 1592 -102
rect 1610 -184 1614 -111
rect 1632 -186 1636 -120
rect 1654 -185 1658 -129
rect 1676 -185 1680 -138
rect 1698 -186 1702 -147
rect 2232 -152 2236 1312
rect 2241 873 2245 1312
rect 2249 876 2253 1312
rect 2281 875 2285 1312
rect 1804 -187 1808 -156
rect 2289 -161 2293 1312
rect 2297 1284 2301 1312
rect 2297 874 2301 1280
rect 2308 56 2309 60
rect 1811 -186 1815 -165
rect 2313 -170 2317 1312
rect 2377 1293 2381 1311
rect 2377 875 2381 1289
rect 2457 920 2461 1314
rect 2497 920 2501 1314
rect 2600 1302 2664 1343
rect 2600 1192 2664 1298
rect 2600 1082 2664 1188
rect 2600 972 2664 1078
rect 2600 862 2664 968
rect 2553 762 2557 811
rect 2600 752 2664 858
rect 2553 652 2557 701
rect 2600 642 2664 748
rect 2553 542 2557 591
rect 2600 532 2664 638
rect 2553 432 2557 481
rect 2600 422 2664 528
rect 2553 322 2557 371
rect 2553 317 2557 318
rect 2600 312 2664 418
rect 2553 212 2557 261
rect 2553 207 2557 208
rect 2600 202 2664 308
rect 2553 102 2557 153
rect 2600 92 2664 198
rect 2385 -80 2389 3
rect 2393 -89 2397 2
rect 2409 -98 2413 -1
rect 2409 -103 2413 -102
rect 2464 -107 2468 2
rect 2520 -116 2524 1
rect 2544 -125 2548 0
rect 2553 -9 2557 41
rect 2560 -134 2564 -2
rect 2574 -143 2578 1
rect 1818 -185 1822 -174
rect 2600 -252 2664 88
rect 2600 -263 2664 -259
rect 2672 1212 2736 1343
rect 2672 1102 2736 1208
rect 2672 992 2736 1098
rect 2672 882 2736 988
rect 2672 772 2736 878
rect 2672 662 2736 768
rect 2672 552 2736 658
rect 2672 442 2736 548
rect 2672 332 2736 438
rect 2672 222 2736 328
rect 2672 112 2736 218
rect 2672 2 2736 108
rect 2672 -277 2736 -2
rect 2672 -289 2736 -284
rect -68 -478 -4 -370
rect -68 -489 -4 -482
<< m3contact >>
rect 16 1238 20 1242
rect 24 1218 28 1222
rect 8 1198 12 1202
rect 136 1238 140 1242
rect 136 958 140 962
rect 88 948 92 952
rect 64 848 68 852
rect 40 828 44 832
rect 0 808 4 812
rect 32 798 36 802
rect 64 738 68 742
rect 40 718 44 722
rect 0 698 4 702
rect 32 688 36 692
rect 64 628 68 632
rect 40 608 44 612
rect 0 588 4 592
rect 32 578 36 582
rect 64 518 68 522
rect 40 498 44 502
rect 0 478 4 482
rect 32 468 36 472
rect 64 408 68 412
rect 40 388 44 392
rect 0 368 4 372
rect 32 358 36 362
rect 64 298 68 302
rect 40 278 44 282
rect 0 258 4 262
rect 392 1278 396 1282
rect 408 1178 412 1182
rect 400 1168 404 1172
rect 400 1158 404 1162
rect 392 1128 396 1132
rect 384 1068 388 1072
rect 376 1048 380 1052
rect 368 1018 372 1022
rect 320 958 324 962
rect 272 948 276 952
rect 248 848 252 852
rect 248 738 252 742
rect 248 628 252 632
rect 248 518 252 522
rect 248 408 252 412
rect 248 298 252 302
rect 32 248 36 252
rect 64 188 68 192
rect 248 188 252 192
rect 40 168 44 172
rect 0 148 4 152
rect 408 1058 412 1062
rect 32 138 36 142
rect 64 78 68 82
rect 248 78 252 82
rect 40 58 44 62
rect 0 38 4 42
rect 552 1258 556 1262
rect 504 958 508 962
rect 456 948 460 952
rect 432 848 436 852
rect 432 738 436 742
rect 432 628 436 632
rect 560 1148 564 1152
rect 432 518 436 522
rect 568 1038 572 1042
rect 432 408 436 412
rect 616 1218 620 1222
rect 664 958 668 962
rect 616 948 620 952
rect 696 938 700 942
rect 592 848 596 852
rect 696 828 700 832
rect 592 738 596 742
rect 617 718 621 722
rect 592 628 596 632
rect 592 518 596 522
rect 592 408 596 412
rect 432 298 436 302
rect 592 298 596 302
rect 432 188 436 192
rect 592 188 596 192
rect 432 78 436 82
rect 592 78 596 82
rect 32 28 36 32
rect 544 -156 548 -152
rect 704 828 708 832
rect 704 718 708 722
rect 704 608 708 612
rect 704 498 708 502
rect 704 388 708 392
rect 704 278 708 282
rect 704 168 708 172
rect 704 58 708 62
rect 768 1258 772 1262
rect 768 1148 772 1152
rect 768 1038 772 1042
rect 800 1278 804 1282
rect 1496 1289 1500 1293
rect 800 1168 804 1172
rect 800 1058 804 1062
rect 816 958 820 962
rect 768 948 772 952
rect 872 938 876 942
rect 768 848 772 852
rect 912 818 916 822
rect 904 808 908 812
rect 768 738 772 742
rect 912 708 916 712
rect 904 698 908 702
rect 768 628 772 632
rect 912 598 916 602
rect 904 588 908 592
rect 768 518 772 522
rect 912 488 916 492
rect 904 478 908 482
rect 768 408 772 412
rect 912 378 916 382
rect 904 368 908 372
rect 768 298 772 302
rect 912 268 916 272
rect 904 258 908 262
rect 768 188 772 192
rect 912 158 916 162
rect 904 148 908 152
rect 768 78 772 82
rect 912 48 916 52
rect 904 38 908 42
rect 1478 -12 1482 -8
rect 1398 -21 1402 -17
rect 1318 -30 1322 -26
rect 1238 -39 1242 -35
rect 1158 -48 1162 -44
rect 1078 -57 1082 -53
rect 696 -165 700 -161
rect 998 -66 1002 -62
rect 617 -174 621 -170
rect 1190 -75 1194 -71
rect 1584 1280 1588 1284
rect 1552 958 1556 962
rect 1504 948 1508 952
rect 1504 778 1508 782
rect 1504 668 1508 672
rect 1504 558 1508 562
rect 1504 448 1508 452
rect 1504 338 1508 342
rect 1504 228 1508 232
rect 1504 118 1508 122
rect 1504 8 1508 12
rect 1760 958 1764 962
rect 1712 948 1716 952
rect 1912 958 1916 962
rect 1864 948 1868 952
rect 2080 1198 2084 1202
rect 2144 958 2148 962
rect 2096 948 2100 952
rect 1848 847 1852 851
rect 2186 848 2190 852
rect 1592 838 1596 842
rect 1616 838 1620 842
rect 1696 838 1700 842
rect 1656 828 1660 832
rect 1672 828 1676 832
rect 2168 838 2172 842
rect 2016 828 2020 832
rect 1840 798 1844 802
rect 1712 788 1716 792
rect 1952 808 1956 812
rect 1976 808 1980 812
rect 1864 778 1868 782
rect 1968 778 1972 782
rect 1592 728 1596 732
rect 1616 728 1620 732
rect 1656 718 1660 722
rect 2176 838 2180 842
rect 2176 826 2180 830
rect 2186 813 2190 817
rect 2176 798 2180 802
rect 2176 778 2180 782
rect 2176 758 2180 762
rect 1688 748 1692 752
rect 2168 748 2172 752
rect 1672 718 1676 722
rect 1592 618 1596 622
rect 1616 618 1620 622
rect 1656 608 1660 612
rect 1672 608 1676 612
rect 1592 508 1596 512
rect 1616 508 1620 512
rect 1656 498 1660 502
rect 1672 498 1676 502
rect 1592 398 1596 402
rect 1616 398 1620 402
rect 1656 388 1660 392
rect 1672 388 1676 392
rect 1592 288 1596 292
rect 1616 288 1620 292
rect 1656 278 1660 282
rect 1672 278 1676 282
rect 1592 178 1596 182
rect 1616 178 1620 182
rect 1656 168 1660 172
rect 1592 68 1596 72
rect 1616 68 1620 72
rect 1656 58 1660 62
rect 1672 168 1676 172
rect 1672 58 1676 62
rect 1529 -2 1533 2
rect 1584 -2 1588 2
rect 1496 -187 1500 -183
rect 1505 -187 1509 -183
rect 1848 737 1852 741
rect 2186 738 2190 742
rect 1696 728 1700 732
rect 2168 728 2172 732
rect 2016 718 2020 722
rect 1840 688 1844 692
rect 1712 678 1716 682
rect 1952 698 1956 702
rect 1976 698 1980 702
rect 1864 668 1868 672
rect 1968 668 1972 672
rect 2176 728 2180 732
rect 2176 716 2180 720
rect 2186 703 2190 707
rect 2176 688 2180 692
rect 2176 668 2180 672
rect 2176 648 2180 652
rect 1704 638 1708 642
rect 2168 638 2172 642
rect 1696 618 1700 622
rect 1696 508 1700 512
rect 1696 398 1700 402
rect 1696 288 1700 292
rect 1696 178 1700 182
rect 1696 68 1700 72
rect 1688 -12 1692 -8
rect 1848 627 1852 631
rect 2186 628 2190 632
rect 2168 618 2172 622
rect 2016 608 2020 612
rect 1840 578 1844 582
rect 1712 568 1716 572
rect 1952 588 1956 592
rect 1976 588 1980 592
rect 1864 558 1868 562
rect 1968 558 1972 562
rect 2176 618 2180 622
rect 2176 606 2180 610
rect 2186 593 2190 597
rect 2176 578 2180 582
rect 2176 558 2180 562
rect 2176 538 2180 542
rect 1792 528 1796 532
rect 2168 528 2172 532
rect 1712 458 1716 462
rect 1712 348 1716 352
rect 1712 238 1716 242
rect 1712 128 1716 132
rect 1712 18 1716 22
rect 1704 -21 1708 -17
rect 1848 517 1852 521
rect 2186 518 2190 522
rect 2168 508 2172 512
rect 2016 498 2020 502
rect 1840 468 1844 472
rect 1952 478 1956 482
rect 1976 478 1980 482
rect 1864 448 1868 452
rect 1968 448 1972 452
rect 2176 508 2180 512
rect 2176 496 2180 500
rect 2186 483 2190 487
rect 2176 468 2180 472
rect 2176 448 2180 452
rect 2176 428 2180 432
rect 1856 418 1860 422
rect 2168 418 2172 422
rect 1848 407 1852 411
rect 1840 358 1844 362
rect 1848 297 1852 301
rect 1840 248 1844 252
rect 1848 187 1852 191
rect 1840 138 1844 142
rect 1848 77 1852 81
rect 1840 28 1844 32
rect 1792 -30 1796 -26
rect 2168 398 2172 402
rect 2016 388 2020 392
rect 1952 368 1956 372
rect 1976 368 1980 372
rect 1864 338 1868 342
rect 1968 338 1972 342
rect 2176 398 2180 402
rect 2176 386 2180 390
rect 2186 373 2190 377
rect 2176 358 2180 362
rect 2176 338 2180 342
rect 2176 318 2180 322
rect 1944 308 1948 312
rect 2168 308 2172 312
rect 1864 228 1868 232
rect 1864 118 1868 122
rect 1864 8 1868 12
rect 1856 -39 1860 -35
rect 2185 298 2189 302
rect 2168 288 2172 292
rect 2016 278 2020 282
rect 1952 258 1956 262
rect 1976 258 1980 262
rect 1968 228 1972 232
rect 2176 288 2180 292
rect 2176 276 2180 280
rect 2185 263 2189 267
rect 2176 248 2180 252
rect 2176 228 2180 232
rect 2176 208 2180 212
rect 1992 198 1996 202
rect 2168 198 2172 202
rect 1952 148 1956 152
rect 1976 148 1980 152
rect 1968 118 1972 122
rect 1952 38 1956 42
rect 1976 38 1980 42
rect 1968 8 1972 12
rect 1944 -48 1948 -44
rect 2186 188 2190 192
rect 2168 178 2172 182
rect 2016 168 2020 172
rect 2024 88 2028 92
rect 2176 178 2180 182
rect 2176 168 2180 172
rect 2186 155 2190 159
rect 2176 138 2180 142
rect 2176 118 2180 122
rect 2176 98 2180 102
rect 2168 88 2172 92
rect 2016 58 2020 62
rect 1992 -57 1996 -53
rect 2186 78 2190 82
rect 2024 -66 2028 -62
rect 2168 68 2172 72
rect 2176 68 2180 72
rect 2176 56 2180 60
rect 2186 43 2190 47
rect 2176 28 2180 32
rect 2176 8 2180 12
rect 2176 -13 2180 -9
rect 2168 -75 2172 -71
rect 1544 -84 1548 -80
rect 1566 -93 1570 -89
rect 1588 -102 1592 -98
rect 1610 -111 1614 -107
rect 1632 -120 1636 -116
rect 1654 -129 1658 -125
rect 1676 -138 1680 -134
rect 1698 -147 1702 -143
rect 1804 -156 1808 -152
rect 2232 -156 2236 -152
rect 2297 1280 2301 1284
rect 1811 -165 1815 -161
rect 2289 -165 2293 -161
rect 2377 1289 2381 1293
rect 2553 758 2557 762
rect 2553 648 2557 652
rect 2553 538 2557 542
rect 2553 428 2557 432
rect 2553 318 2557 322
rect 2553 208 2557 212
rect 2553 98 2557 102
rect 2385 -84 2389 -80
rect 2393 -93 2397 -89
rect 2409 -102 2413 -98
rect 2464 -111 2468 -107
rect 2520 -120 2524 -116
rect 2553 -13 2557 -9
rect 2544 -129 2548 -125
rect 2560 -138 2564 -134
rect 2574 -147 2578 -143
rect 1818 -174 1822 -170
rect 2313 -174 2317 -170
<< metal3 >>
rect 1495 1293 2382 1294
rect 1495 1289 1496 1293
rect 1500 1289 2377 1293
rect 2381 1289 2382 1293
rect 1495 1288 2382 1289
rect 1583 1284 2302 1285
rect 391 1282 805 1283
rect 391 1278 392 1282
rect 396 1278 800 1282
rect 804 1278 805 1282
rect 1583 1280 1584 1284
rect 1588 1280 2297 1284
rect 2301 1280 2302 1284
rect 1583 1279 2302 1280
rect 391 1277 805 1278
rect 551 1262 773 1263
rect 551 1258 552 1262
rect 556 1258 768 1262
rect 772 1258 773 1262
rect 551 1257 773 1258
rect 15 1242 141 1243
rect 15 1238 16 1242
rect 20 1238 136 1242
rect 140 1238 141 1242
rect 15 1237 141 1238
rect 23 1222 956 1223
rect 23 1218 24 1222
rect 28 1218 616 1222
rect 620 1218 956 1222
rect 23 1217 956 1218
rect 7 1202 2085 1203
rect 7 1198 8 1202
rect 12 1198 2080 1202
rect 2084 1198 2085 1202
rect 7 1197 2085 1198
rect 407 1182 892 1183
rect 407 1178 408 1182
rect 412 1178 892 1182
rect 407 1177 892 1178
rect 399 1172 805 1173
rect 399 1168 400 1172
rect 404 1168 800 1172
rect 804 1168 805 1172
rect 399 1167 805 1168
rect 399 1162 860 1163
rect 399 1158 400 1162
rect 404 1158 860 1162
rect 399 1157 860 1158
rect 559 1152 773 1153
rect 559 1148 560 1152
rect 564 1148 768 1152
rect 772 1148 773 1152
rect 559 1147 773 1148
rect 391 1132 828 1133
rect 391 1128 392 1132
rect 396 1128 828 1132
rect 391 1127 828 1128
rect 383 1072 892 1073
rect 383 1068 384 1072
rect 388 1068 892 1072
rect 383 1067 892 1068
rect 407 1062 805 1063
rect 407 1058 408 1062
rect 412 1058 800 1062
rect 804 1058 805 1062
rect 407 1057 805 1058
rect 375 1052 860 1053
rect 375 1048 376 1052
rect 380 1048 860 1052
rect 375 1047 860 1048
rect 567 1042 773 1043
rect 567 1038 568 1042
rect 572 1038 768 1042
rect 772 1038 773 1042
rect 567 1037 773 1038
rect 367 1022 828 1023
rect 367 1018 368 1022
rect 372 1018 828 1022
rect 367 1017 828 1018
rect 135 962 2149 963
rect 135 958 136 962
rect 140 958 320 962
rect 324 958 504 962
rect 508 958 664 962
rect 668 958 816 962
rect 820 958 1552 962
rect 1556 958 1760 962
rect 1764 958 1912 962
rect 1916 958 2144 962
rect 2148 958 2149 962
rect 135 957 2149 958
rect 87 952 2101 953
rect 87 948 88 952
rect 92 948 272 952
rect 276 948 456 952
rect 460 948 616 952
rect 620 948 768 952
rect 772 948 1504 952
rect 1508 948 1712 952
rect 1716 948 1864 952
rect 1868 948 2096 952
rect 2100 948 2101 952
rect 87 947 2101 948
rect 695 942 877 943
rect 695 938 696 942
rect 700 938 872 942
rect 876 938 877 942
rect 695 937 877 938
rect -17 852 773 853
rect -17 848 64 852
rect 68 848 248 852
rect 252 848 432 852
rect 436 848 592 852
rect 596 848 768 852
rect 772 848 773 852
rect -17 847 773 848
rect 1847 852 2191 853
rect 1847 851 2186 852
rect 1847 847 1848 851
rect 1852 848 2186 851
rect 2190 848 2191 852
rect 1852 847 2191 848
rect 1847 846 1853 847
rect -17 842 1621 843
rect -17 838 1592 842
rect 1596 838 1616 842
rect 1620 838 1621 842
rect -17 837 1621 838
rect 1695 842 2182 843
rect 1695 838 1696 842
rect 1700 838 2168 842
rect 2172 838 2176 842
rect 2180 838 2182 842
rect 1695 837 2182 838
rect -17 832 45 833
rect -17 828 40 832
rect 44 828 45 832
rect -17 827 45 828
rect 695 832 1661 833
rect 695 828 696 832
rect 700 828 704 832
rect 708 828 1656 832
rect 1660 828 1661 832
rect 695 827 1661 828
rect 1671 832 2021 833
rect 1671 828 1672 832
rect 1676 828 2016 832
rect 2020 828 2021 832
rect 1671 827 2021 828
rect 2175 830 2198 831
rect 2175 826 2176 830
rect 2180 826 2198 830
rect 2175 825 2198 826
rect 911 822 925 823
rect 911 818 912 822
rect 916 818 925 822
rect 911 817 925 818
rect 2185 817 2198 818
rect 2185 813 2186 817
rect 2190 813 2198 817
rect -1 812 1981 813
rect 2185 812 2198 813
rect -1 808 0 812
rect 4 808 904 812
rect 908 808 1952 812
rect 1956 808 1976 812
rect 1980 808 1981 812
rect -1 807 1981 808
rect 31 802 2181 803
rect 31 798 32 802
rect 36 798 1840 802
rect 1844 798 2176 802
rect 2180 798 2181 802
rect 31 797 2181 798
rect 1487 792 1717 793
rect 1487 788 1712 792
rect 1716 788 1717 792
rect 1487 787 1717 788
rect 1487 782 1509 783
rect 1487 778 1504 782
rect 1508 778 1509 782
rect 1487 777 1509 778
rect 1863 782 2182 783
rect 1863 778 1864 782
rect 1868 778 1968 782
rect 1972 778 2176 782
rect 2180 778 2182 782
rect 1863 777 2182 778
rect 2175 762 2558 763
rect 2175 758 2176 762
rect 2180 758 2553 762
rect 2557 758 2558 762
rect 2175 757 2558 758
rect 1687 752 2173 753
rect 1687 748 1688 752
rect 1692 748 2168 752
rect 2172 748 2173 752
rect 1687 747 2173 748
rect -17 742 773 743
rect -17 738 64 742
rect 68 738 248 742
rect 252 738 432 742
rect 436 738 592 742
rect 596 738 768 742
rect 772 738 773 742
rect -17 737 773 738
rect 1847 742 2191 743
rect 1847 741 2186 742
rect 1847 737 1848 741
rect 1852 738 2186 741
rect 2190 738 2191 742
rect 1852 737 2191 738
rect 1847 736 1853 737
rect -17 732 1621 733
rect -17 728 1592 732
rect 1596 728 1616 732
rect 1620 728 1621 732
rect -17 727 1621 728
rect 1695 732 2182 733
rect 1695 728 1696 732
rect 1700 728 2168 732
rect 2172 728 2176 732
rect 2180 728 2182 732
rect 1695 727 2182 728
rect -17 722 45 723
rect -17 718 40 722
rect 44 718 45 722
rect -17 717 45 718
rect 615 722 1661 723
rect 615 718 617 722
rect 621 718 704 722
rect 708 718 1656 722
rect 1660 718 1661 722
rect 615 717 1661 718
rect 1671 722 2021 723
rect 1671 718 1672 722
rect 1676 718 2016 722
rect 2020 718 2021 722
rect 1671 717 2021 718
rect 2175 720 2198 721
rect 2175 716 2176 720
rect 2180 716 2198 720
rect 2175 715 2198 716
rect 911 712 925 713
rect 911 708 912 712
rect 916 708 925 712
rect 911 707 925 708
rect 2185 707 2198 708
rect 2185 703 2186 707
rect 2190 703 2198 707
rect -1 702 1981 703
rect 2185 702 2198 703
rect -1 698 0 702
rect 4 698 904 702
rect 908 698 1952 702
rect 1956 698 1976 702
rect 1980 698 1981 702
rect -1 697 1981 698
rect 31 692 2181 693
rect 31 688 32 692
rect 36 688 1840 692
rect 1844 688 2176 692
rect 2180 688 2181 692
rect 31 687 2181 688
rect 1487 682 1717 683
rect 1487 678 1712 682
rect 1716 678 1717 682
rect 1487 677 1717 678
rect 1487 672 1509 673
rect 1487 668 1504 672
rect 1508 668 1509 672
rect 1487 667 1509 668
rect 1863 672 2182 673
rect 1863 668 1864 672
rect 1868 668 1968 672
rect 1972 668 2176 672
rect 2180 668 2182 672
rect 1863 667 2182 668
rect 2175 652 2558 653
rect 2175 648 2176 652
rect 2180 648 2553 652
rect 2557 648 2558 652
rect 2175 647 2558 648
rect 1703 642 2173 643
rect 1703 638 1704 642
rect 1708 638 2168 642
rect 2172 638 2173 642
rect 1703 637 2173 638
rect -17 632 773 633
rect -17 628 64 632
rect 68 628 248 632
rect 252 628 432 632
rect 436 628 592 632
rect 596 628 768 632
rect 772 628 773 632
rect -17 627 773 628
rect 1847 632 2191 633
rect 1847 631 2186 632
rect 1847 627 1848 631
rect 1852 628 2186 631
rect 2190 628 2191 632
rect 1852 627 2191 628
rect 1847 626 1853 627
rect -17 622 1621 623
rect -17 618 1592 622
rect 1596 618 1616 622
rect 1620 618 1621 622
rect -17 617 1621 618
rect 1695 622 2182 623
rect 1695 618 1696 622
rect 1700 618 2168 622
rect 2172 618 2176 622
rect 2180 618 2182 622
rect 1695 617 2182 618
rect -17 612 45 613
rect -17 608 40 612
rect 44 608 45 612
rect -17 607 45 608
rect 703 612 1661 613
rect 703 608 704 612
rect 708 608 1656 612
rect 1660 608 1661 612
rect 703 607 1661 608
rect 1671 612 2021 613
rect 1671 608 1672 612
rect 1676 608 2016 612
rect 2020 608 2021 612
rect 1671 607 2021 608
rect 2175 610 2198 611
rect 2175 606 2176 610
rect 2180 606 2198 610
rect 2175 605 2198 606
rect 911 602 925 603
rect 911 598 912 602
rect 916 598 925 602
rect 911 597 925 598
rect 2185 597 2198 598
rect 2185 593 2186 597
rect 2190 593 2198 597
rect -1 592 1981 593
rect 2185 592 2198 593
rect -1 588 0 592
rect 4 588 904 592
rect 908 588 1952 592
rect 1956 588 1976 592
rect 1980 588 1981 592
rect -1 587 1981 588
rect 31 582 2181 583
rect 31 578 32 582
rect 36 578 1840 582
rect 1844 578 2176 582
rect 2180 578 2181 582
rect 31 577 2181 578
rect 1487 572 1717 573
rect 1487 568 1712 572
rect 1716 568 1717 572
rect 1487 567 1717 568
rect 1487 562 1509 563
rect 1487 558 1504 562
rect 1508 558 1509 562
rect 1487 557 1509 558
rect 1863 562 2182 563
rect 1863 558 1864 562
rect 1868 558 1968 562
rect 1972 558 2176 562
rect 2180 558 2182 562
rect 1863 557 2182 558
rect 2175 542 2558 543
rect 2175 538 2176 542
rect 2180 538 2553 542
rect 2557 538 2558 542
rect 2175 537 2558 538
rect 1791 532 2173 533
rect 1791 528 1792 532
rect 1796 528 2168 532
rect 2172 528 2173 532
rect 1791 527 2173 528
rect -17 522 773 523
rect -17 518 64 522
rect 68 518 248 522
rect 252 518 432 522
rect 436 518 592 522
rect 596 518 768 522
rect 772 518 773 522
rect -17 517 773 518
rect 1847 522 2191 523
rect 1847 521 2186 522
rect 1847 517 1848 521
rect 1852 518 2186 521
rect 2190 518 2191 522
rect 1852 517 2191 518
rect 1847 516 1853 517
rect -17 512 1621 513
rect -17 508 1592 512
rect 1596 508 1616 512
rect 1620 508 1621 512
rect -17 507 1621 508
rect 1695 512 2182 513
rect 1695 508 1696 512
rect 1700 508 2168 512
rect 2172 508 2176 512
rect 2180 508 2182 512
rect 1695 507 2182 508
rect -17 502 45 503
rect -17 498 40 502
rect 44 498 45 502
rect -17 497 45 498
rect 703 502 1661 503
rect 703 498 704 502
rect 708 498 1656 502
rect 1660 498 1661 502
rect 703 497 1661 498
rect 1671 502 2021 503
rect 1671 498 1672 502
rect 1676 498 2016 502
rect 2020 498 2021 502
rect 1671 497 2021 498
rect 2175 500 2198 501
rect 2175 496 2176 500
rect 2180 496 2198 500
rect 2175 495 2198 496
rect 911 492 925 493
rect 911 488 912 492
rect 916 488 925 492
rect 911 487 925 488
rect 2185 487 2198 488
rect 2185 483 2186 487
rect 2190 483 2198 487
rect -1 482 1981 483
rect 2185 482 2198 483
rect -1 478 0 482
rect 4 478 904 482
rect 908 478 1952 482
rect 1956 478 1976 482
rect 1980 478 1981 482
rect -1 477 1981 478
rect 31 472 2181 473
rect 31 468 32 472
rect 36 468 1840 472
rect 1844 468 2176 472
rect 2180 468 2181 472
rect 31 467 2181 468
rect 1487 462 1717 463
rect 1487 458 1712 462
rect 1716 458 1717 462
rect 1487 457 1717 458
rect 1487 452 1509 453
rect 1487 448 1504 452
rect 1508 448 1509 452
rect 1487 447 1509 448
rect 1863 452 2182 453
rect 1863 448 1864 452
rect 1868 448 1968 452
rect 1972 448 2176 452
rect 2180 448 2182 452
rect 1863 447 2182 448
rect 2175 432 2558 433
rect 2175 428 2176 432
rect 2180 428 2553 432
rect 2557 428 2558 432
rect 2175 427 2558 428
rect 1855 422 2173 423
rect 1855 418 1856 422
rect 1860 418 2168 422
rect 2172 418 2173 422
rect 1855 417 2173 418
rect -17 412 773 413
rect -17 408 64 412
rect 68 408 248 412
rect 252 408 432 412
rect 436 408 592 412
rect 596 408 768 412
rect 772 408 773 412
rect -17 407 773 408
rect 1847 411 2191 413
rect 1847 407 1848 411
rect 1852 407 2191 411
rect 1847 406 1853 407
rect -17 402 1621 403
rect -17 398 1592 402
rect 1596 398 1616 402
rect 1620 398 1621 402
rect -17 397 1621 398
rect 1695 402 2182 403
rect 1695 398 1696 402
rect 1700 398 2168 402
rect 2172 398 2176 402
rect 2180 398 2182 402
rect 1695 397 2182 398
rect -17 392 45 393
rect -17 388 40 392
rect 44 388 45 392
rect -17 387 45 388
rect 703 392 1661 393
rect 703 388 704 392
rect 708 388 1656 392
rect 1660 388 1661 392
rect 703 387 1661 388
rect 1671 392 2021 393
rect 1671 388 1672 392
rect 1676 388 2016 392
rect 2020 388 2021 392
rect 1671 387 2021 388
rect 2175 390 2198 391
rect 2175 386 2176 390
rect 2180 386 2198 390
rect 2175 385 2198 386
rect 911 382 925 383
rect 911 378 912 382
rect 916 378 925 382
rect 911 377 925 378
rect 2185 377 2198 378
rect 2185 373 2186 377
rect 2190 373 2198 377
rect -1 372 1981 373
rect 2185 372 2198 373
rect -1 368 0 372
rect 4 368 904 372
rect 908 368 1952 372
rect 1956 368 1976 372
rect 1980 368 1981 372
rect -1 367 1981 368
rect 31 362 2181 363
rect 31 358 32 362
rect 36 358 1840 362
rect 1844 358 2176 362
rect 2180 358 2181 362
rect 31 357 2181 358
rect 1487 352 1717 353
rect 1487 348 1712 352
rect 1716 348 1717 352
rect 1487 347 1717 348
rect 1487 342 1509 343
rect 1487 338 1504 342
rect 1508 338 1509 342
rect 1487 337 1509 338
rect 1863 342 2182 343
rect 1863 338 1864 342
rect 1868 338 1968 342
rect 1972 338 2176 342
rect 2180 338 2182 342
rect 1863 337 2182 338
rect 2175 322 2558 323
rect 2175 318 2176 322
rect 2180 318 2553 322
rect 2557 318 2558 322
rect 2175 317 2558 318
rect 1943 312 2173 313
rect 1943 308 1944 312
rect 1948 308 2168 312
rect 2172 308 2173 312
rect 1943 307 2173 308
rect -17 302 773 303
rect -17 298 64 302
rect 68 298 248 302
rect 252 298 432 302
rect 436 298 592 302
rect 596 298 768 302
rect 772 298 773 302
rect -17 297 773 298
rect 1847 302 2190 303
rect 1847 301 2185 302
rect 1847 297 1848 301
rect 1852 298 2185 301
rect 2189 298 2190 302
rect 1852 297 2190 298
rect 1847 296 1853 297
rect -17 292 1621 293
rect -17 288 1592 292
rect 1596 288 1616 292
rect 1620 288 1621 292
rect -17 287 1621 288
rect 1695 292 2182 293
rect 1695 288 1696 292
rect 1700 288 2168 292
rect 2172 288 2176 292
rect 2180 288 2182 292
rect 1695 287 2182 288
rect -17 282 45 283
rect -17 278 40 282
rect 44 278 45 282
rect -17 277 45 278
rect 703 282 1661 283
rect 703 278 704 282
rect 708 278 1656 282
rect 1660 278 1661 282
rect 703 277 1661 278
rect 1671 282 2021 283
rect 1671 278 1672 282
rect 1676 278 2016 282
rect 2020 278 2021 282
rect 1671 277 2021 278
rect 2175 280 2198 281
rect 2175 276 2176 280
rect 2180 276 2198 280
rect 2175 275 2198 276
rect 911 272 925 273
rect 911 268 912 272
rect 916 268 925 272
rect 911 267 925 268
rect 2184 267 2198 268
rect 2184 263 2185 267
rect 2189 263 2198 267
rect -1 262 1981 263
rect 2184 262 2198 263
rect -1 258 0 262
rect 4 258 904 262
rect 908 258 1952 262
rect 1956 258 1976 262
rect 1980 258 1981 262
rect -1 257 1981 258
rect 31 252 2181 253
rect 31 248 32 252
rect 36 248 1840 252
rect 1844 248 2176 252
rect 2180 248 2181 252
rect 31 247 2181 248
rect 1487 242 1717 243
rect 1487 238 1712 242
rect 1716 238 1717 242
rect 1487 237 1717 238
rect 1487 232 1509 233
rect 1487 228 1504 232
rect 1508 228 1509 232
rect 1487 227 1509 228
rect 1863 232 2182 233
rect 1863 228 1864 232
rect 1868 228 1968 232
rect 1972 228 2176 232
rect 2180 228 2182 232
rect 1863 227 2182 228
rect 2175 212 2558 213
rect 2175 208 2176 212
rect 2180 208 2553 212
rect 2557 208 2558 212
rect 2175 207 2558 208
rect 1991 202 2173 203
rect 1991 198 1992 202
rect 1996 198 2168 202
rect 2172 198 2173 202
rect 1991 197 2173 198
rect -17 192 773 193
rect -17 188 64 192
rect 68 188 248 192
rect 252 188 432 192
rect 436 188 592 192
rect 596 188 768 192
rect 772 188 773 192
rect -17 187 773 188
rect 1847 192 2191 193
rect 1847 191 2186 192
rect 1847 187 1848 191
rect 1852 188 2186 191
rect 2190 188 2191 192
rect 1852 187 2191 188
rect 1847 186 1853 187
rect -17 182 1621 183
rect -17 178 1592 182
rect 1596 178 1616 182
rect 1620 178 1621 182
rect -17 177 1621 178
rect 1695 182 2182 183
rect 1695 178 1696 182
rect 1700 178 2168 182
rect 2172 178 2176 182
rect 2180 178 2182 182
rect 1695 177 2182 178
rect -17 172 45 173
rect -17 168 40 172
rect 44 168 45 172
rect -17 167 45 168
rect 703 172 1661 173
rect 703 168 704 172
rect 708 168 1656 172
rect 1660 168 1661 172
rect 703 167 1661 168
rect 1671 172 2021 173
rect 1671 168 1672 172
rect 1676 168 2016 172
rect 2020 168 2021 172
rect 1671 167 2021 168
rect 2175 172 2198 173
rect 2175 168 2176 172
rect 2180 168 2198 172
rect 2175 167 2198 168
rect 911 162 925 163
rect 911 158 912 162
rect 916 158 925 162
rect 911 157 925 158
rect 2185 159 2198 160
rect 2185 155 2186 159
rect 2190 155 2198 159
rect 2185 154 2198 155
rect -1 152 1981 153
rect -1 148 0 152
rect 4 148 904 152
rect 908 148 1952 152
rect 1956 148 1976 152
rect 1980 148 1981 152
rect -1 147 1981 148
rect 31 142 2181 143
rect 31 138 32 142
rect 36 138 1840 142
rect 1844 138 2176 142
rect 2180 138 2181 142
rect 31 137 2181 138
rect 1487 132 1717 133
rect 1487 128 1712 132
rect 1716 128 1717 132
rect 1487 127 1717 128
rect 1487 122 1509 123
rect 1487 118 1504 122
rect 1508 118 1509 122
rect 1487 117 1509 118
rect 1863 122 2182 123
rect 1863 118 1864 122
rect 1868 118 1968 122
rect 1972 118 2176 122
rect 2180 118 2182 122
rect 1863 117 2182 118
rect 2175 102 2558 103
rect 2175 98 2176 102
rect 2180 98 2553 102
rect 2557 98 2558 102
rect 2175 97 2558 98
rect 2023 92 2173 93
rect 2023 88 2024 92
rect 2028 88 2168 92
rect 2172 88 2173 92
rect 2023 87 2173 88
rect -17 82 773 83
rect -17 78 64 82
rect 68 78 248 82
rect 252 78 432 82
rect 436 78 592 82
rect 596 78 768 82
rect 772 78 773 82
rect -17 77 773 78
rect 1847 82 2191 83
rect 1847 81 2186 82
rect 1847 77 1848 81
rect 1852 78 2186 81
rect 2190 78 2191 82
rect 1852 77 2191 78
rect 1847 76 1853 77
rect -17 72 1621 73
rect -17 68 1592 72
rect 1596 68 1616 72
rect 1620 68 1621 72
rect -17 67 1621 68
rect 1695 72 2182 73
rect 1695 68 1696 72
rect 1700 68 2168 72
rect 2172 68 2176 72
rect 2180 68 2182 72
rect 1695 67 2182 68
rect -17 62 45 63
rect -17 58 40 62
rect 44 58 45 62
rect -17 57 45 58
rect 703 62 1661 63
rect 703 58 704 62
rect 708 58 1656 62
rect 1660 58 1661 62
rect 703 57 1661 58
rect 1671 62 2021 63
rect 1671 58 1672 62
rect 1676 58 2016 62
rect 2020 58 2021 62
rect 1671 57 2021 58
rect 2175 60 2198 61
rect 2175 56 2176 60
rect 2180 56 2198 60
rect 2175 55 2198 56
rect 911 52 925 53
rect 911 48 912 52
rect 916 48 925 52
rect 911 47 925 48
rect 2185 47 2197 48
rect 2185 43 2186 47
rect 2190 43 2197 47
rect -1 42 1981 43
rect 2185 42 2197 43
rect -1 38 0 42
rect 4 38 904 42
rect 908 38 1952 42
rect 1956 38 1976 42
rect 1980 38 1981 42
rect -1 37 1981 38
rect 31 32 2181 33
rect 31 28 32 32
rect 36 28 1840 32
rect 1844 28 2176 32
rect 2180 28 2181 32
rect 31 27 2181 28
rect 1487 22 1717 23
rect 1487 18 1712 22
rect 1716 18 1717 22
rect 1487 17 1717 18
rect 1487 12 1509 13
rect 1487 8 1504 12
rect 1508 8 1509 12
rect 1487 7 1509 8
rect 1863 12 2182 13
rect 1863 8 1864 12
rect 1868 8 1968 12
rect 1972 8 2176 12
rect 2180 8 2182 12
rect 1863 7 2182 8
rect 1528 2 1589 3
rect 1528 -2 1529 2
rect 1533 -2 1584 2
rect 1588 -2 1589 2
rect 1528 -3 1589 -2
rect 1477 -8 1693 -7
rect 1477 -12 1478 -8
rect 1482 -12 1688 -8
rect 1692 -12 1693 -8
rect 1477 -13 1693 -12
rect 2175 -9 2558 -8
rect 2175 -13 2176 -9
rect 2180 -13 2553 -9
rect 2557 -13 2558 -9
rect 2175 -14 2558 -13
rect 1397 -17 1709 -16
rect 1397 -21 1398 -17
rect 1402 -21 1704 -17
rect 1708 -21 1709 -17
rect 1397 -22 1709 -21
rect 1317 -26 1797 -25
rect 1317 -30 1318 -26
rect 1322 -30 1792 -26
rect 1796 -30 1797 -26
rect 1317 -31 1797 -30
rect 1237 -35 1861 -34
rect 1237 -39 1238 -35
rect 1242 -39 1856 -35
rect 1860 -39 1861 -35
rect 1237 -40 1861 -39
rect 1157 -44 1949 -43
rect 1157 -48 1158 -44
rect 1162 -48 1944 -44
rect 1948 -48 1949 -44
rect 1157 -49 1949 -48
rect 1077 -53 1997 -52
rect 1077 -57 1078 -53
rect 1082 -57 1992 -53
rect 1996 -57 1997 -53
rect 1077 -58 1997 -57
rect 997 -62 2029 -61
rect 997 -66 998 -62
rect 1002 -66 2024 -62
rect 2028 -66 2029 -62
rect 997 -67 2029 -66
rect 1189 -71 2173 -70
rect 1189 -75 1190 -71
rect 1194 -75 2168 -71
rect 2172 -75 2173 -71
rect 1189 -76 2173 -75
rect 1543 -80 2390 -79
rect 1543 -84 1544 -80
rect 1548 -84 2385 -80
rect 2389 -84 2390 -80
rect 1543 -85 2390 -84
rect 1565 -89 2398 -88
rect 1565 -93 1566 -89
rect 1570 -93 2393 -89
rect 2397 -93 2398 -89
rect 1565 -94 2398 -93
rect 1587 -98 2414 -97
rect 1587 -102 1588 -98
rect 1592 -102 2409 -98
rect 2413 -102 2414 -98
rect 1587 -103 2414 -102
rect 1609 -107 2469 -106
rect 1609 -111 1610 -107
rect 1614 -111 2464 -107
rect 2468 -111 2469 -107
rect 1609 -112 2469 -111
rect 1631 -116 2525 -115
rect 1631 -120 1632 -116
rect 1636 -120 2520 -116
rect 2524 -120 2525 -116
rect 1631 -121 2525 -120
rect 1653 -125 2549 -124
rect 1653 -129 1654 -125
rect 1658 -129 2544 -125
rect 2548 -129 2549 -125
rect 1653 -130 2549 -129
rect 1675 -134 2565 -133
rect 1675 -138 1676 -134
rect 1680 -138 2560 -134
rect 2564 -138 2565 -134
rect 1675 -139 2565 -138
rect 1697 -143 2579 -142
rect 1697 -147 1698 -143
rect 1702 -147 2574 -143
rect 2578 -147 2579 -143
rect 1697 -148 2579 -147
rect 543 -152 2237 -151
rect 543 -156 544 -152
rect 548 -156 1804 -152
rect 1808 -156 2232 -152
rect 2236 -156 2237 -152
rect 543 -157 2237 -156
rect 695 -161 2294 -160
rect 695 -165 696 -161
rect 700 -165 1811 -161
rect 1815 -165 2289 -161
rect 2293 -165 2294 -161
rect 695 -166 2294 -165
rect 616 -170 2318 -169
rect 616 -174 617 -170
rect 621 -174 1818 -170
rect 1822 -174 2313 -170
rect 2317 -174 2318 -170
rect 616 -175 2318 -174
rect 1495 -183 1510 -182
rect 1495 -187 1496 -183
rect 1500 -187 1505 -183
rect 1509 -187 1510 -183
rect 1495 -188 1510 -187
use mux2_c_1x  mux2_c_1x_0
timestamp 1484534138
transform 1 0 760 0 1 1210
box -6 -4 66 96
use mux2_c_1x  mux2_c_1x_1
timestamp 1484534138
transform 1 0 760 0 1 1100
box -6 -4 66 96
use mux2_c_1x  mux2_c_1x_2
timestamp 1484534138
transform 1 0 760 0 1 990
box -6 -4 66 96
use mux2_1x_8  mux2_1x_8_0
timestamp 1484532969
transform 1 0 0 0 1 0
box -6 -4 50 976
use flopen_1x_8  flopen_1x_8_0
timestamp 1484532171
transform 1 0 48 0 1 0
box -6 -4 138 976
use flopen_1x_8  flopen_1x_8_1
timestamp 1484532171
transform 1 0 232 0 1 0
box -6 -4 138 976
use flopen_1x_8  flopen_1x_8_2
timestamp 1484532171
transform 1 0 416 0 1 0
box -6 -4 138 976
use flopen_1x_8  flopen_1x_8_3
timestamp 1484532171
transform 1 0 576 0 1 0
box -6 -4 138 976
use flop_1x_8  flop_1x_8_0
timestamp 1484532171
transform 1 0 761 0 1 0
box -7 -4 105 976
use mux2_1x_8  mux2_1x_8_1
timestamp 1484532969
transform 1 0 872 0 1 0
box -6 -4 50 976
use flop_1x_8  flop_1x_8_1
timestamp 1484532171
transform 1 0 1497 0 1 0
box -7 -4 105 976
use mux4_1x_8  mux4_1x_8_0
timestamp 1484532969
transform 1 0 1600 0 1 0
box -6 -4 106 976
use flop_1x_8  flop_1x_8_2
timestamp 1484532171
transform 1 0 1705 0 1 0
box -7 -4 105 976
use mux2_1x_8  mux2_1x_8_2
timestamp 1484532969
transform 1 0 1808 0 1 0
box -6 -4 50 976
use flop_1x_8  flop_1x_8_3
timestamp 1484532171
transform 1 0 1857 0 1 0
box -7 -4 105 976
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 1960 0 1 0
box -6 -4 82 976
use flopenr_1x_8  flopenr_1x_8_0
timestamp 1484532171
transform 1 0 2040 0 1 0
box -6 -4 147 976
use alt_alu_8  alt_alu_8_0
timestamp 1493690245
transform 1 0 2187 0 1 -4
box 0 0 410 982
use regramarray_dp  regramarray_dp_0
timestamp 1488938149
transform 1 0 920 0 1 0
box -102 -5 578 1306
use array_sh_sg  array_sh_sg_0
timestamp 1493690245
transform 1 0 944 0 1 -484
box 0 -64 1539 301
<< labels >>
rlabel metal2 697 -14 697 -14 1 shamt1
rlabel metal2 2291 1310 2291 1310 1 k1
rlabel metal2 545 -6 545 -6 1 shamt2
rlabel metal2 2708 1340 2708 1340 5 Gnd!
rlabel metal2 2625 1340 2625 1340 5 Vdd!
rlabel metal2 1480 -116 1480 -116 1 sc7
rlabel metal2 1400 -119 1400 -119 1 sc6
rlabel metal2 1320 -117 1320 -117 1 sc5
rlabel metal2 1240 -117 1240 -117 1 sc4
rlabel metal2 1191 -120 1191 -120 1 sc0
rlabel metal2 1160 -119 1160 -119 1 sc3
rlabel metal2 1080 -123 1080 -123 1 sc2
rlabel metal2 1000 -122 1000 -122 1 sc1
rlabel metal2 1700 -183 1700 -183 1 y0
rlabel metal2 1678 -183 1678 -183 1 y1
rlabel metal2 1656 -184 1656 -184 1 y2
rlabel metal2 1634 -184 1634 -184 1 y3
rlabel metal2 1611 -183 1611 -183 1 y4
rlabel metal2 1590 -183 1590 -183 1 y5
rlabel metal2 1568 -183 1568 -183 1 y6
rlabel metal2 1546 -183 1546 -183 1 y7
rlabel m3contact 2178 120 2178 120 1 result1
rlabel m3contact 2178 230 2178 230 1 result2
rlabel m3contact 2178 340 2178 340 1 result3
rlabel m3contact 2178 450 2178 450 1 result4
rlabel m3contact 2178 560 2178 560 1 result5
rlabel m3contact 2178 670 2178 670 1 result6
rlabel m3contact 2178 780 2178 780 1 result7
rlabel metal2 2315 1310 2315 1310 1 k0
rlabel m3contact 2178 10 2178 10 1 result0
rlabel metal2 2499 1312 2499 1312 1 op1
rlabel metal2 2459 1312 2459 1312 1 op0
rlabel metal2 2379 1309 2379 1309 1 op2
rlabel metal2 2299 1310 2299 1310 1 op3
rlabel metal2 2283 1310 2283 1310 1 op4
rlabel metal2 2251 1310 2251 1310 1 op5
rlabel metal2 2243 1310 2243 1310 1 op6
rlabel metal3 2195 814 2195 814 1 a7
rlabel metal3 2194 704 2194 704 1 a6
rlabel metal3 2195 595 2195 595 1 a5
rlabel metal3 2195 484 2195 484 1 a4
rlabel metal3 2195 374 2195 374 1 a3
rlabel metal3 2196 264 2196 264 1 a2
rlabel metal3 2195 156 2195 156 1 a1
rlabel metal3 2195 44 2195 44 1 a0
rlabel metal2 2234 1310 2234 1310 1 k2
rlabel metal2 1498 1310 1498 1310 1 arith
rlabel metal2 1586 1310 1586 1310 1 right
rlabel metal2 1690 -6 1690 -6 1 b7
rlabel metal2 1706 -5 1706 -5 1 b6
rlabel metal2 1794 -5 1794 -5 1 b5
rlabel metal2 1858 -5 1858 -5 1 b4
rlabel metal2 1946 -6 1946 -6 1 b3
rlabel metal2 1994 -5 1994 -5 1 b2
rlabel metal2 2026 -5 2026 -5 1 b1
rlabel metal2 2170 -11 2170 -11 1 b0
rlabel metal3 2180 10 2180 10 1 result0
rlabel metal3 2180 70 2180 70 1 b0
rlabel metal3 2180 80 2180 80 1 a0
rlabel metal2 -34 1336 -34 1336 1 Gnd!
rlabel metal2 -106 1336 -106 1336 1 Vdd!
rlabel metal3 -15 60 -15 60 1 adr0
rlabel metal3 -15 70 -15 70 1 writedata0
rlabel metal3 -14 80 -14 80 1 memdata0
rlabel metal3 -15 170 -15 170 1 adr1
rlabel metal3 -15 180 -15 180 1 writedata1
rlabel metal3 -14 190 -14 190 1 memdata1
rlabel metal3 -14 280 -14 280 1 adr2
rlabel metal3 -14 290 -14 290 1 writedata2
rlabel metal3 -13 300 -13 300 1 memdata2
rlabel metal3 -14 390 -14 390 1 adr3
rlabel metal3 -13 400 -13 400 1 writedata3
rlabel metal3 -14 409 -14 409 1 memdata3
rlabel metal3 -14 500 -14 500 1 adr4
rlabel metal3 -14 510 -14 510 1 writedata4
rlabel metal3 -14 519 -14 519 1 memdata4
rlabel metal3 -15 610 -15 610 1 adr5
rlabel metal3 -15 619 -15 619 1 writedata5
rlabel metal3 -14 630 -14 630 1 memdata5
rlabel metal3 -14 721 -14 721 1 adr6
rlabel metal3 -15 729 -15 729 1 writedata6
rlabel metal3 -15 739 -15 739 1 memdata6
rlabel metal3 -13 831 -13 831 1 adr7
rlabel metal3 -13 839 -13 839 1 writedata7
rlabel metal3 -13 850 -13 850 1 memdata7
rlabel metal2 26 1310 26 1310 1 ph2
rlabel metal2 18 1310 18 1310 1 ph1
rlabel metal2 10 1310 10 1310 1 reset
rlabel metal2 2 1310 2 1310 1 iord
rlabel metal2 58 1310 58 1310 1 irwrite_3_
rlabel metal2 186 1309 186 1309 1 op_5_
rlabel metal2 194 1310 194 1310 1 op_4_
rlabel metal2 202 1309 202 1309 1 op_3_
rlabel metal2 210 1311 210 1311 1 op_2_
rlabel metal2 218 1308 218 1308 1 op_1_
rlabel metal2 226 1310 226 1310 1 op_0_
rlabel metal2 242 1310 242 1310 1 irwrite_2_
rlabel metal2 426 1310 426 1310 1 irwrite_1_
rlabel metal2 586 1310 586 1310 1 irwrite_0_
rlabel metal2 698 1310 698 1310 1 memtoreg
rlabel metal2 714 1309 714 1309 1 funct_5_
rlabel metal2 722 1310 722 1310 1 funct_4_
rlabel metal2 730 1309 730 1309 1 funct_3_
rlabel metal2 738 1311 738 1311 1 funct_2_
rlabel metal2 746 1308 746 1308 1 funct_1_
rlabel metal2 753 1309 753 1309 1 funct_0_
rlabel metal2 794 1309 794 1309 1 regdst
rlabel metal2 961 1310 961 1310 1 regwrite
rlabel metal2 1601 1310 1601 1310 1 alusrcb_0_
rlabel metal2 1633 1310 1633 1310 1 alusrcb_1_
rlabel metal2 1809 1309 1809 1309 1 alusrca
rlabel metal2 1962 1309 1962 1309 1 pcsrc_0
rlabel metal2 1994 1310 1994 1310 1 pcsrc_1_
rlabel metal2 2050 1309 2050 1309 1 pcen
rlabel metal2 619 -10 619 -10 1 shamt0
<< end >>
