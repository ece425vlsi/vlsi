magic
tech scmos
timestamp 1493737109
<< m2contact >>
rect -7 -7 7 7
<< end >>
