magic
tech scmos
timestamp 1488306180
<< m2contact >>
rect -2 -2 2 2
<< end >>
