magic
tech scmos
timestamp 1399650201
<< metal1 >>
rect 2 -1 3 -0
rect 3 -1 4 -0
rect 4 -1 5 -0
rect 5 -1 6 -0
rect 6 -1 7 -0
rect 7 -1 8 -0
rect 8 -1 9 -0
rect 9 -1 10 -0
rect 10 -1 11 -0
rect 11 -1 12 -0
rect 12 -1 13 -0
rect 13 -1 14 -0
rect 14 -1 15 -0
rect 15 -1 16 -0
rect 16 -1 17 -0
rect 17 -1 18 -0
rect 18 -1 19 -0
rect 19 -1 20 -0
rect 20 -1 21 -0
rect 21 -1 22 -0
rect 22 -1 23 -0
rect 23 -1 24 -0
rect 24 -1 25 -0
rect 25 -1 26 -0
rect 26 -1 27 -0
rect 27 -1 28 -0
rect 28 -1 29 -0
rect 29 -1 30 -0
rect 30 -1 31 -0
rect 31 -1 32 -0
rect 32 -1 33 -0
rect 33 -1 34 -0
rect 34 -1 35 -0
rect 35 -1 36 -0
rect 36 -1 37 -0
rect 37 -1 38 -0
rect 38 -1 39 -0
rect 39 -1 40 -0
rect 40 -1 41 -0
rect 41 -1 42 -0
rect 42 -1 43 -0
rect 43 -1 44 -0
rect 44 -1 45 -0
rect 45 -1 46 -0
rect 46 -1 47 -0
rect 47 -1 48 -0
rect 48 -1 49 -0
rect 49 -1 50 -0
rect 50 -1 51 -0
rect 51 -1 52 -0
rect 52 -1 53 -0
rect 53 -1 54 -0
rect 54 -1 55 -0
rect 55 -1 56 -0
rect 56 -1 57 -0
rect 57 -1 58 -0
rect 58 -1 59 -0
rect 59 -1 60 -0
rect 60 -1 61 -0
rect 61 -1 62 -0
rect 62 -1 63 -0
rect 63 -1 64 -0
rect 64 -1 65 -0
rect 65 -1 66 -0
rect 66 -1 67 -0
rect 67 -1 68 -0
rect 68 -1 69 -0
rect 69 -1 70 -0
rect 70 -1 71 -0
rect 71 -1 72 -0
rect 72 -1 73 -0
rect 73 -1 74 -0
rect 74 -1 75 -0
rect 75 -1 76 -0
rect 76 -1 77 -0
rect 77 -1 78 -0
rect 78 -1 79 -0
rect 79 -1 80 -0
rect 80 -1 81 -0
rect 81 -1 82 -0
rect 82 -1 83 -0
rect 83 -1 84 -0
rect 84 -1 85 -0
rect 85 -1 86 -0
rect 86 -1 87 -0
rect 87 -1 88 -0
rect 88 -1 89 -0
rect 89 -1 90 -0
rect 90 -1 91 -0
rect 91 -1 92 -0
rect 92 -1 93 -0
rect 93 -1 94 -0
rect 94 -1 95 -0
rect 95 -1 96 -0
rect 96 -1 97 -0
rect 97 -1 98 -0
rect 98 -1 99 -0
rect 99 -1 100 -0
rect 100 -1 101 -0
rect 101 -1 102 -0
rect 102 -1 103 -0
rect 103 -1 104 -0
rect 104 -1 105 -0
rect 105 -1 106 -0
rect 106 -1 107 -0
rect 107 -1 108 -0
rect 108 -1 109 -0
rect 109 -1 110 -0
rect 110 -1 111 -0
rect 111 -1 112 -0
rect 112 -1 113 -0
rect 113 -1 114 -0
rect 114 -1 115 -0
rect 115 -1 116 -0
rect 116 -1 117 -0
rect 117 -1 118 -0
rect 118 -1 119 -0
rect 119 -1 120 -0
rect 120 -1 121 -0
rect 121 -1 122 -0
rect 122 -1 123 -0
rect 123 -1 124 -0
rect 124 -1 125 -0
rect 125 -1 126 -0
rect 126 -1 127 -0
rect 127 -1 128 -0
rect 128 -1 129 -0
rect 129 -1 130 -0
rect 130 -1 131 -0
rect 131 -1 132 -0
rect 132 -1 133 -0
rect 133 -1 134 -0
rect 134 -1 135 -0
rect 135 -1 136 -0
rect 136 -1 137 -0
rect 137 -1 138 -0
rect 138 -1 139 -0
rect 139 -1 140 -0
rect 140 -1 141 -0
rect 141 -1 142 -0
rect 142 -1 143 -0
rect 143 -1 144 -0
rect 144 -1 145 -0
rect 145 -1 146 -0
rect 146 -1 147 -0
rect 147 -1 148 -0
rect 148 -1 149 -0
rect 149 -1 150 -0
rect 150 -1 151 -0
rect 151 -1 152 -0
rect 152 -1 153 -0
rect 153 -1 154 -0
rect 154 -1 155 -0
rect 155 -1 156 -0
rect 156 -1 157 -0
rect 157 -1 158 -0
rect 158 -1 159 -0
rect 159 -1 160 -0
rect 160 -1 161 -0
rect 161 -1 162 -0
rect 162 -1 163 -0
rect 163 -1 164 -0
rect 164 -1 165 -0
rect 165 -1 166 -0
rect 166 -1 167 -0
rect 167 -1 168 -0
rect 168 -1 169 -0
rect 169 -1 170 -0
rect 170 -1 171 -0
rect 171 -1 172 -0
rect 172 -1 173 -0
rect 173 -1 174 -0
rect 174 -1 175 -0
rect 175 -1 176 -0
rect 176 -1 177 -0
rect 177 -1 178 -0
rect 178 -1 179 -0
rect 179 -1 180 -0
rect 180 -1 181 -0
rect 181 -1 182 -0
rect 182 -1 183 -0
rect 183 -1 184 -0
rect 184 -1 185 -0
rect 185 -1 186 -0
rect 186 -1 187 -0
rect 187 -1 188 -0
rect 188 -1 189 -0
rect 189 -1 190 -0
rect 190 -1 191 -0
rect 191 -1 192 -0
rect 192 -1 193 -0
rect 193 -1 194 -0
rect 194 -1 195 -0
rect 195 -1 196 -0
rect 196 -1 197 -0
rect 197 -1 198 -0
rect 198 -1 199 -0
rect 199 -1 200 -0
rect 200 -1 201 -0
rect 201 -1 202 -0
rect 202 -1 203 -0
rect 203 -1 204 -0
rect 204 -1 205 -0
rect 205 -1 206 -0
rect 206 -1 207 -0
rect 207 -1 208 -0
rect 208 -1 209 -0
rect 209 -1 210 -0
rect 210 -1 211 -0
rect 211 -1 212 -0
rect 212 -1 213 -0
rect 213 -1 214 -0
rect 214 -1 215 -0
rect 215 -1 216 -0
rect 216 -1 217 -0
rect 217 -1 218 -0
rect 218 -1 219 -0
rect 219 -1 220 -0
rect 220 -1 221 -0
rect 221 -1 222 -0
rect 222 -1 223 -0
rect 223 -1 224 -0
rect 224 -1 225 -0
rect 225 -1 226 -0
rect 226 -1 227 -0
rect 227 -1 228 -0
rect 228 -1 229 -0
rect 229 -1 230 -0
rect 230 -1 231 -0
rect 231 -1 232 -0
rect 232 -1 233 -0
rect 233 -1 234 -0
rect 234 -1 235 -0
rect 235 -1 236 -0
rect 236 -1 237 -0
rect 237 -1 238 -0
rect 238 -1 239 -0
rect 239 -1 240 -0
rect 240 -1 241 -0
rect 241 -1 242 -0
rect 242 -1 243 -0
rect 243 -1 244 -0
rect 244 -1 245 -0
rect 245 -1 246 -0
rect 246 -1 247 -0
rect 247 -1 248 -0
rect 248 -1 249 -0
rect 249 -1 250 -0
rect 250 -1 251 -0
rect 251 -1 252 -0
rect 252 -1 253 -0
rect 253 -1 254 -0
rect 254 -1 255 -0
rect 255 -1 256 -0
rect 256 -1 257 -0
rect 257 -1 258 -0
rect 258 -1 259 -0
rect 259 -1 260 -0
rect 260 -1 261 -0
rect 261 -1 262 -0
rect 262 -1 263 -0
rect 263 -1 264 -0
rect 264 -1 265 -0
rect 265 -1 266 -0
rect 266 -1 267 -0
rect 267 -1 268 -0
rect 268 -1 269 -0
rect 269 -1 270 -0
rect 270 -1 271 -0
rect 271 -1 272 -0
rect 272 -1 273 -0
rect 273 -1 274 -0
rect 274 -1 275 -0
rect 275 -1 276 -0
rect 276 -1 277 -0
rect 277 -1 278 -0
rect 278 -1 279 -0
rect 279 -1 280 -0
rect 280 -1 281 -0
rect 281 -1 282 -0
rect 282 -1 283 -0
rect 283 -1 284 -0
rect 284 -1 285 -0
rect 285 -1 286 -0
rect 286 -1 287 -0
rect 287 -1 288 -0
rect 288 -1 289 -0
rect 289 -1 290 -0
rect 290 -1 291 -0
rect 291 -1 292 -0
rect 292 -1 293 -0
rect 293 -1 294 -0
rect 294 -1 295 -0
rect 295 -1 296 -0
rect 296 -1 297 -0
rect 297 -1 298 -0
rect 298 -1 299 -0
rect 299 -1 300 -0
rect 300 -1 301 -0
rect 301 -1 302 -0
rect 302 -1 303 -0
rect 303 -1 304 -0
rect 304 -1 305 -0
rect 305 -1 306 -0
rect 306 -1 307 -0
rect 307 -1 308 -0
rect 308 -1 309 -0
rect 309 -1 310 -0
rect 310 -1 311 -0
rect 311 -1 312 -0
rect 312 -1 313 -0
rect 313 -1 314 -0
rect 314 -1 315 -0
rect 315 -1 316 -0
rect 316 -1 317 -0
rect 317 -1 318 -0
rect 318 -1 319 -0
rect 319 -1 320 -0
rect 320 -1 321 -0
rect 321 -1 322 -0
rect 322 -1 323 -0
rect 323 -1 324 -0
rect 324 -1 325 -0
rect 325 -1 326 -0
rect 326 -1 327 -0
rect 327 -1 328 -0
rect 328 -1 329 -0
rect 329 -1 330 -0
rect 330 -1 331 -0
rect 331 -1 332 -0
rect 332 -1 333 -0
rect 333 -1 334 -0
rect 334 -1 335 -0
rect 335 -1 336 -0
rect 336 -1 337 -0
rect 337 -1 338 -0
rect 338 -1 339 -0
rect 339 -1 340 -0
rect 340 -1 341 -0
rect 341 -1 342 -0
rect 342 -1 343 -0
rect 343 -1 344 -0
rect 344 -1 345 -0
rect 345 -1 346 -0
rect 346 -1 347 -0
rect 347 -1 348 -0
rect 348 -1 349 -0
rect 349 -1 350 -0
rect 350 -1 351 -0
rect 351 -1 352 -0
rect 352 -1 353 -0
rect 353 -1 354 -0
rect 354 -1 355 -0
rect 355 -1 356 -0
rect 356 -1 357 -0
rect 357 -1 358 -0
rect 358 -1 359 -0
rect 359 -1 360 -0
rect 360 -1 361 -0
rect 361 -1 362 -0
rect 362 -1 363 -0
rect 363 -1 364 -0
rect 364 -1 365 -0
rect 365 -1 366 -0
rect 366 -1 367 -0
rect 367 -1 368 -0
rect 368 -1 369 -0
rect 369 -1 370 -0
rect 370 -1 371 -0
rect 371 -1 372 -0
rect 372 -1 373 -0
rect 373 -1 374 -0
rect 374 -1 375 -0
rect 375 -1 376 -0
rect 376 -1 377 -0
rect 377 -1 378 -0
rect 378 -1 379 -0
rect 379 -1 380 -0
rect 380 -1 381 -0
rect 381 -1 382 -0
rect 382 -1 383 -0
rect 383 -1 384 -0
rect 384 -1 385 -0
rect 385 -1 386 -0
rect 386 -1 387 -0
rect 387 -1 388 -0
rect 388 -1 389 -0
rect 389 -1 390 -0
rect 390 -1 391 -0
rect 391 -1 392 -0
rect 392 -1 393 -0
rect 393 -1 394 -0
rect 394 -1 395 -0
rect 395 -1 396 -0
rect 396 -1 397 -0
rect 397 -1 398 -0
rect 398 -1 399 -0
rect 399 -1 400 -0
rect 400 -1 401 -0
rect 401 -1 402 -0
rect 402 -1 403 -0
rect 403 -1 404 -0
rect 404 -1 405 -0
rect 405 -1 406 -0
rect 406 -1 407 -0
rect 407 -1 408 -0
rect 408 -1 409 -0
rect 409 -1 410 -0
rect 410 -1 411 -0
rect 411 -1 412 -0
rect 412 -1 413 -0
rect 413 -1 414 -0
rect 414 -1 415 -0
rect 415 -1 416 -0
rect 416 -1 417 -0
rect 417 -1 418 -0
rect 418 -1 419 -0
rect 419 -1 420 -0
rect 420 -1 421 -0
rect 421 -1 422 -0
rect 422 -1 423 -0
rect 423 -1 424 -0
rect 424 -1 425 -0
rect 425 -1 426 -0
rect 426 -1 427 -0
rect 427 -1 428 -0
rect 428 -1 429 -0
rect 429 -1 430 -0
rect 430 -1 431 -0
rect 431 -1 432 -0
rect 432 -1 433 -0
rect 433 -1 434 -0
rect 434 -1 435 -0
rect 435 -1 436 -0
rect 436 -1 437 -0
rect 437 -1 438 -0
rect 438 -1 439 -0
rect 439 -1 440 -0
rect 440 -1 441 -0
rect 441 -1 442 -0
rect 442 -1 443 -0
rect 443 -1 444 -0
rect 444 -1 445 -0
rect 445 -1 446 -0
rect 446 -1 447 -0
rect 447 -1 448 -0
rect 448 -1 449 -0
rect 449 -1 450 -0
rect 450 -1 451 -0
rect 451 -1 452 -0
rect 452 -1 453 -0
rect 453 -1 454 -0
rect 454 -1 455 -0
rect 455 -1 456 -0
rect 456 -1 457 -0
rect 457 -1 458 -0
rect 458 -1 459 -0
rect 459 -1 460 -0
rect 460 -1 461 -0
rect 461 -1 462 -0
rect 462 -1 463 -0
rect 463 -1 464 -0
rect 464 -1 465 -0
rect 465 -1 466 -0
rect 466 -1 467 -0
rect 467 -1 468 -0
rect 468 -1 469 -0
rect 469 -1 470 -0
rect 470 -1 471 -0
rect 471 -1 472 -0
rect 472 -1 473 -0
rect 473 -1 474 -0
rect 474 -1 475 -0
rect 475 -1 476 -0
rect 476 -1 477 -0
rect 477 -1 478 -0
rect 478 -1 479 -0
rect 479 -1 480 -0
rect 2 -2 3 -1
rect 3 -2 4 -1
rect 4 -2 5 -1
rect 5 -2 6 -1
rect 6 -2 7 -1
rect 7 -2 8 -1
rect 8 -2 9 -1
rect 9 -2 10 -1
rect 10 -2 11 -1
rect 11 -2 12 -1
rect 12 -2 13 -1
rect 13 -2 14 -1
rect 14 -2 15 -1
rect 15 -2 16 -1
rect 16 -2 17 -1
rect 17 -2 18 -1
rect 18 -2 19 -1
rect 19 -2 20 -1
rect 20 -2 21 -1
rect 21 -2 22 -1
rect 22 -2 23 -1
rect 23 -2 24 -1
rect 24 -2 25 -1
rect 25 -2 26 -1
rect 26 -2 27 -1
rect 27 -2 28 -1
rect 28 -2 29 -1
rect 29 -2 30 -1
rect 30 -2 31 -1
rect 31 -2 32 -1
rect 32 -2 33 -1
rect 33 -2 34 -1
rect 34 -2 35 -1
rect 35 -2 36 -1
rect 36 -2 37 -1
rect 37 -2 38 -1
rect 38 -2 39 -1
rect 39 -2 40 -1
rect 40 -2 41 -1
rect 41 -2 42 -1
rect 42 -2 43 -1
rect 43 -2 44 -1
rect 44 -2 45 -1
rect 45 -2 46 -1
rect 46 -2 47 -1
rect 47 -2 48 -1
rect 48 -2 49 -1
rect 49 -2 50 -1
rect 50 -2 51 -1
rect 51 -2 52 -1
rect 52 -2 53 -1
rect 53 -2 54 -1
rect 54 -2 55 -1
rect 55 -2 56 -1
rect 56 -2 57 -1
rect 57 -2 58 -1
rect 58 -2 59 -1
rect 59 -2 60 -1
rect 60 -2 61 -1
rect 61 -2 62 -1
rect 62 -2 63 -1
rect 63 -2 64 -1
rect 64 -2 65 -1
rect 65 -2 66 -1
rect 66 -2 67 -1
rect 67 -2 68 -1
rect 68 -2 69 -1
rect 69 -2 70 -1
rect 70 -2 71 -1
rect 71 -2 72 -1
rect 72 -2 73 -1
rect 73 -2 74 -1
rect 74 -2 75 -1
rect 75 -2 76 -1
rect 76 -2 77 -1
rect 77 -2 78 -1
rect 78 -2 79 -1
rect 79 -2 80 -1
rect 80 -2 81 -1
rect 81 -2 82 -1
rect 82 -2 83 -1
rect 83 -2 84 -1
rect 84 -2 85 -1
rect 85 -2 86 -1
rect 86 -2 87 -1
rect 87 -2 88 -1
rect 88 -2 89 -1
rect 89 -2 90 -1
rect 90 -2 91 -1
rect 91 -2 92 -1
rect 92 -2 93 -1
rect 93 -2 94 -1
rect 94 -2 95 -1
rect 95 -2 96 -1
rect 96 -2 97 -1
rect 97 -2 98 -1
rect 98 -2 99 -1
rect 99 -2 100 -1
rect 100 -2 101 -1
rect 101 -2 102 -1
rect 102 -2 103 -1
rect 103 -2 104 -1
rect 104 -2 105 -1
rect 105 -2 106 -1
rect 106 -2 107 -1
rect 107 -2 108 -1
rect 108 -2 109 -1
rect 109 -2 110 -1
rect 110 -2 111 -1
rect 111 -2 112 -1
rect 112 -2 113 -1
rect 113 -2 114 -1
rect 114 -2 115 -1
rect 115 -2 116 -1
rect 116 -2 117 -1
rect 117 -2 118 -1
rect 118 -2 119 -1
rect 119 -2 120 -1
rect 120 -2 121 -1
rect 121 -2 122 -1
rect 122 -2 123 -1
rect 123 -2 124 -1
rect 124 -2 125 -1
rect 125 -2 126 -1
rect 126 -2 127 -1
rect 127 -2 128 -1
rect 128 -2 129 -1
rect 129 -2 130 -1
rect 130 -2 131 -1
rect 131 -2 132 -1
rect 132 -2 133 -1
rect 133 -2 134 -1
rect 134 -2 135 -1
rect 135 -2 136 -1
rect 136 -2 137 -1
rect 137 -2 138 -1
rect 138 -2 139 -1
rect 139 -2 140 -1
rect 140 -2 141 -1
rect 141 -2 142 -1
rect 142 -2 143 -1
rect 143 -2 144 -1
rect 144 -2 145 -1
rect 145 -2 146 -1
rect 146 -2 147 -1
rect 147 -2 148 -1
rect 148 -2 149 -1
rect 149 -2 150 -1
rect 150 -2 151 -1
rect 151 -2 152 -1
rect 152 -2 153 -1
rect 153 -2 154 -1
rect 154 -2 155 -1
rect 155 -2 156 -1
rect 156 -2 157 -1
rect 157 -2 158 -1
rect 158 -2 159 -1
rect 159 -2 160 -1
rect 160 -2 161 -1
rect 161 -2 162 -1
rect 162 -2 163 -1
rect 163 -2 164 -1
rect 164 -2 165 -1
rect 165 -2 166 -1
rect 166 -2 167 -1
rect 167 -2 168 -1
rect 168 -2 169 -1
rect 169 -2 170 -1
rect 170 -2 171 -1
rect 171 -2 172 -1
rect 172 -2 173 -1
rect 173 -2 174 -1
rect 174 -2 175 -1
rect 175 -2 176 -1
rect 176 -2 177 -1
rect 177 -2 178 -1
rect 178 -2 179 -1
rect 179 -2 180 -1
rect 180 -2 181 -1
rect 181 -2 182 -1
rect 182 -2 183 -1
rect 183 -2 184 -1
rect 184 -2 185 -1
rect 185 -2 186 -1
rect 186 -2 187 -1
rect 187 -2 188 -1
rect 188 -2 189 -1
rect 189 -2 190 -1
rect 190 -2 191 -1
rect 191 -2 192 -1
rect 192 -2 193 -1
rect 193 -2 194 -1
rect 194 -2 195 -1
rect 195 -2 196 -1
rect 196 -2 197 -1
rect 197 -2 198 -1
rect 198 -2 199 -1
rect 199 -2 200 -1
rect 200 -2 201 -1
rect 201 -2 202 -1
rect 202 -2 203 -1
rect 203 -2 204 -1
rect 204 -2 205 -1
rect 205 -2 206 -1
rect 206 -2 207 -1
rect 207 -2 208 -1
rect 208 -2 209 -1
rect 209 -2 210 -1
rect 210 -2 211 -1
rect 211 -2 212 -1
rect 212 -2 213 -1
rect 213 -2 214 -1
rect 214 -2 215 -1
rect 215 -2 216 -1
rect 216 -2 217 -1
rect 217 -2 218 -1
rect 218 -2 219 -1
rect 219 -2 220 -1
rect 220 -2 221 -1
rect 221 -2 222 -1
rect 222 -2 223 -1
rect 223 -2 224 -1
rect 224 -2 225 -1
rect 225 -2 226 -1
rect 226 -2 227 -1
rect 227 -2 228 -1
rect 228 -2 229 -1
rect 229 -2 230 -1
rect 230 -2 231 -1
rect 231 -2 232 -1
rect 232 -2 233 -1
rect 233 -2 234 -1
rect 234 -2 235 -1
rect 235 -2 236 -1
rect 236 -2 237 -1
rect 237 -2 238 -1
rect 238 -2 239 -1
rect 239 -2 240 -1
rect 240 -2 241 -1
rect 241 -2 242 -1
rect 242 -2 243 -1
rect 243 -2 244 -1
rect 244 -2 245 -1
rect 245 -2 246 -1
rect 246 -2 247 -1
rect 247 -2 248 -1
rect 248 -2 249 -1
rect 249 -2 250 -1
rect 250 -2 251 -1
rect 251 -2 252 -1
rect 252 -2 253 -1
rect 253 -2 254 -1
rect 254 -2 255 -1
rect 255 -2 256 -1
rect 256 -2 257 -1
rect 257 -2 258 -1
rect 258 -2 259 -1
rect 259 -2 260 -1
rect 260 -2 261 -1
rect 261 -2 262 -1
rect 262 -2 263 -1
rect 263 -2 264 -1
rect 264 -2 265 -1
rect 265 -2 266 -1
rect 266 -2 267 -1
rect 267 -2 268 -1
rect 268 -2 269 -1
rect 269 -2 270 -1
rect 270 -2 271 -1
rect 271 -2 272 -1
rect 272 -2 273 -1
rect 273 -2 274 -1
rect 274 -2 275 -1
rect 275 -2 276 -1
rect 276 -2 277 -1
rect 277 -2 278 -1
rect 278 -2 279 -1
rect 279 -2 280 -1
rect 280 -2 281 -1
rect 281 -2 282 -1
rect 282 -2 283 -1
rect 283 -2 284 -1
rect 284 -2 285 -1
rect 285 -2 286 -1
rect 286 -2 287 -1
rect 287 -2 288 -1
rect 288 -2 289 -1
rect 289 -2 290 -1
rect 290 -2 291 -1
rect 291 -2 292 -1
rect 292 -2 293 -1
rect 293 -2 294 -1
rect 294 -2 295 -1
rect 295 -2 296 -1
rect 296 -2 297 -1
rect 297 -2 298 -1
rect 298 -2 299 -1
rect 299 -2 300 -1
rect 300 -2 301 -1
rect 301 -2 302 -1
rect 302 -2 303 -1
rect 303 -2 304 -1
rect 304 -2 305 -1
rect 305 -2 306 -1
rect 306 -2 307 -1
rect 307 -2 308 -1
rect 308 -2 309 -1
rect 309 -2 310 -1
rect 310 -2 311 -1
rect 311 -2 312 -1
rect 312 -2 313 -1
rect 313 -2 314 -1
rect 314 -2 315 -1
rect 315 -2 316 -1
rect 316 -2 317 -1
rect 317 -2 318 -1
rect 318 -2 319 -1
rect 319 -2 320 -1
rect 320 -2 321 -1
rect 321 -2 322 -1
rect 322 -2 323 -1
rect 323 -2 324 -1
rect 324 -2 325 -1
rect 325 -2 326 -1
rect 326 -2 327 -1
rect 327 -2 328 -1
rect 328 -2 329 -1
rect 329 -2 330 -1
rect 330 -2 331 -1
rect 331 -2 332 -1
rect 332 -2 333 -1
rect 333 -2 334 -1
rect 334 -2 335 -1
rect 335 -2 336 -1
rect 336 -2 337 -1
rect 337 -2 338 -1
rect 338 -2 339 -1
rect 339 -2 340 -1
rect 340 -2 341 -1
rect 341 -2 342 -1
rect 342 -2 343 -1
rect 343 -2 344 -1
rect 344 -2 345 -1
rect 345 -2 346 -1
rect 346 -2 347 -1
rect 347 -2 348 -1
rect 348 -2 349 -1
rect 349 -2 350 -1
rect 350 -2 351 -1
rect 351 -2 352 -1
rect 352 -2 353 -1
rect 353 -2 354 -1
rect 354 -2 355 -1
rect 355 -2 356 -1
rect 356 -2 357 -1
rect 357 -2 358 -1
rect 358 -2 359 -1
rect 359 -2 360 -1
rect 360 -2 361 -1
rect 361 -2 362 -1
rect 362 -2 363 -1
rect 363 -2 364 -1
rect 364 -2 365 -1
rect 365 -2 366 -1
rect 366 -2 367 -1
rect 367 -2 368 -1
rect 368 -2 369 -1
rect 369 -2 370 -1
rect 370 -2 371 -1
rect 371 -2 372 -1
rect 372 -2 373 -1
rect 373 -2 374 -1
rect 374 -2 375 -1
rect 375 -2 376 -1
rect 376 -2 377 -1
rect 377 -2 378 -1
rect 378 -2 379 -1
rect 379 -2 380 -1
rect 380 -2 381 -1
rect 381 -2 382 -1
rect 382 -2 383 -1
rect 383 -2 384 -1
rect 384 -2 385 -1
rect 385 -2 386 -1
rect 386 -2 387 -1
rect 387 -2 388 -1
rect 388 -2 389 -1
rect 389 -2 390 -1
rect 390 -2 391 -1
rect 391 -2 392 -1
rect 392 -2 393 -1
rect 393 -2 394 -1
rect 394 -2 395 -1
rect 395 -2 396 -1
rect 396 -2 397 -1
rect 397 -2 398 -1
rect 398 -2 399 -1
rect 399 -2 400 -1
rect 400 -2 401 -1
rect 401 -2 402 -1
rect 402 -2 403 -1
rect 403 -2 404 -1
rect 404 -2 405 -1
rect 405 -2 406 -1
rect 406 -2 407 -1
rect 407 -2 408 -1
rect 408 -2 409 -1
rect 409 -2 410 -1
rect 410 -2 411 -1
rect 411 -2 412 -1
rect 412 -2 413 -1
rect 413 -2 414 -1
rect 414 -2 415 -1
rect 415 -2 416 -1
rect 416 -2 417 -1
rect 417 -2 418 -1
rect 418 -2 419 -1
rect 419 -2 420 -1
rect 420 -2 421 -1
rect 421 -2 422 -1
rect 422 -2 423 -1
rect 423 -2 424 -1
rect 424 -2 425 -1
rect 425 -2 426 -1
rect 426 -2 427 -1
rect 427 -2 428 -1
rect 428 -2 429 -1
rect 429 -2 430 -1
rect 430 -2 431 -1
rect 431 -2 432 -1
rect 432 -2 433 -1
rect 433 -2 434 -1
rect 434 -2 435 -1
rect 435 -2 436 -1
rect 436 -2 437 -1
rect 437 -2 438 -1
rect 438 -2 439 -1
rect 439 -2 440 -1
rect 440 -2 441 -1
rect 441 -2 442 -1
rect 442 -2 443 -1
rect 443 -2 444 -1
rect 444 -2 445 -1
rect 445 -2 446 -1
rect 446 -2 447 -1
rect 447 -2 448 -1
rect 448 -2 449 -1
rect 449 -2 450 -1
rect 450 -2 451 -1
rect 451 -2 452 -1
rect 452 -2 453 -1
rect 453 -2 454 -1
rect 454 -2 455 -1
rect 455 -2 456 -1
rect 456 -2 457 -1
rect 457 -2 458 -1
rect 458 -2 459 -1
rect 459 -2 460 -1
rect 460 -2 461 -1
rect 461 -2 462 -1
rect 462 -2 463 -1
rect 463 -2 464 -1
rect 464 -2 465 -1
rect 465 -2 466 -1
rect 466 -2 467 -1
rect 467 -2 468 -1
rect 468 -2 469 -1
rect 469 -2 470 -1
rect 470 -2 471 -1
rect 471 -2 472 -1
rect 472 -2 473 -1
rect 473 -2 474 -1
rect 474 -2 475 -1
rect 475 -2 476 -1
rect 476 -2 477 -1
rect 477 -2 478 -1
rect 478 -2 479 -1
rect 479 -2 480 -1
rect 2 -3 3 -2
rect 3 -3 4 -2
rect 4 -3 5 -2
rect 5 -3 6 -2
rect 6 -3 7 -2
rect 7 -3 8 -2
rect 8 -3 9 -2
rect 9 -3 10 -2
rect 10 -3 11 -2
rect 11 -3 12 -2
rect 12 -3 13 -2
rect 13 -3 14 -2
rect 14 -3 15 -2
rect 15 -3 16 -2
rect 16 -3 17 -2
rect 17 -3 18 -2
rect 18 -3 19 -2
rect 19 -3 20 -2
rect 20 -3 21 -2
rect 21 -3 22 -2
rect 22 -3 23 -2
rect 23 -3 24 -2
rect 24 -3 25 -2
rect 25 -3 26 -2
rect 26 -3 27 -2
rect 27 -3 28 -2
rect 28 -3 29 -2
rect 29 -3 30 -2
rect 30 -3 31 -2
rect 31 -3 32 -2
rect 32 -3 33 -2
rect 33 -3 34 -2
rect 34 -3 35 -2
rect 35 -3 36 -2
rect 36 -3 37 -2
rect 37 -3 38 -2
rect 38 -3 39 -2
rect 39 -3 40 -2
rect 40 -3 41 -2
rect 41 -3 42 -2
rect 42 -3 43 -2
rect 43 -3 44 -2
rect 44 -3 45 -2
rect 45 -3 46 -2
rect 46 -3 47 -2
rect 47 -3 48 -2
rect 48 -3 49 -2
rect 49 -3 50 -2
rect 50 -3 51 -2
rect 51 -3 52 -2
rect 52 -3 53 -2
rect 53 -3 54 -2
rect 54 -3 55 -2
rect 55 -3 56 -2
rect 56 -3 57 -2
rect 57 -3 58 -2
rect 58 -3 59 -2
rect 59 -3 60 -2
rect 60 -3 61 -2
rect 61 -3 62 -2
rect 62 -3 63 -2
rect 63 -3 64 -2
rect 64 -3 65 -2
rect 65 -3 66 -2
rect 66 -3 67 -2
rect 67 -3 68 -2
rect 68 -3 69 -2
rect 69 -3 70 -2
rect 70 -3 71 -2
rect 71 -3 72 -2
rect 72 -3 73 -2
rect 73 -3 74 -2
rect 74 -3 75 -2
rect 75 -3 76 -2
rect 76 -3 77 -2
rect 77 -3 78 -2
rect 78 -3 79 -2
rect 79 -3 80 -2
rect 80 -3 81 -2
rect 81 -3 82 -2
rect 82 -3 83 -2
rect 83 -3 84 -2
rect 84 -3 85 -2
rect 85 -3 86 -2
rect 86 -3 87 -2
rect 87 -3 88 -2
rect 88 -3 89 -2
rect 89 -3 90 -2
rect 90 -3 91 -2
rect 91 -3 92 -2
rect 92 -3 93 -2
rect 93 -3 94 -2
rect 94 -3 95 -2
rect 95 -3 96 -2
rect 96 -3 97 -2
rect 97 -3 98 -2
rect 98 -3 99 -2
rect 99 -3 100 -2
rect 100 -3 101 -2
rect 101 -3 102 -2
rect 102 -3 103 -2
rect 103 -3 104 -2
rect 104 -3 105 -2
rect 105 -3 106 -2
rect 106 -3 107 -2
rect 107 -3 108 -2
rect 108 -3 109 -2
rect 109 -3 110 -2
rect 110 -3 111 -2
rect 111 -3 112 -2
rect 112 -3 113 -2
rect 113 -3 114 -2
rect 114 -3 115 -2
rect 115 -3 116 -2
rect 116 -3 117 -2
rect 117 -3 118 -2
rect 118 -3 119 -2
rect 119 -3 120 -2
rect 120 -3 121 -2
rect 121 -3 122 -2
rect 122 -3 123 -2
rect 123 -3 124 -2
rect 124 -3 125 -2
rect 125 -3 126 -2
rect 126 -3 127 -2
rect 127 -3 128 -2
rect 128 -3 129 -2
rect 129 -3 130 -2
rect 130 -3 131 -2
rect 131 -3 132 -2
rect 132 -3 133 -2
rect 133 -3 134 -2
rect 134 -3 135 -2
rect 135 -3 136 -2
rect 136 -3 137 -2
rect 137 -3 138 -2
rect 138 -3 139 -2
rect 139 -3 140 -2
rect 140 -3 141 -2
rect 141 -3 142 -2
rect 142 -3 143 -2
rect 143 -3 144 -2
rect 144 -3 145 -2
rect 145 -3 146 -2
rect 146 -3 147 -2
rect 147 -3 148 -2
rect 148 -3 149 -2
rect 149 -3 150 -2
rect 150 -3 151 -2
rect 151 -3 152 -2
rect 152 -3 153 -2
rect 153 -3 154 -2
rect 154 -3 155 -2
rect 155 -3 156 -2
rect 156 -3 157 -2
rect 157 -3 158 -2
rect 158 -3 159 -2
rect 159 -3 160 -2
rect 160 -3 161 -2
rect 161 -3 162 -2
rect 162 -3 163 -2
rect 163 -3 164 -2
rect 164 -3 165 -2
rect 165 -3 166 -2
rect 166 -3 167 -2
rect 167 -3 168 -2
rect 168 -3 169 -2
rect 169 -3 170 -2
rect 170 -3 171 -2
rect 171 -3 172 -2
rect 172 -3 173 -2
rect 173 -3 174 -2
rect 174 -3 175 -2
rect 175 -3 176 -2
rect 176 -3 177 -2
rect 177 -3 178 -2
rect 178 -3 179 -2
rect 179 -3 180 -2
rect 180 -3 181 -2
rect 181 -3 182 -2
rect 182 -3 183 -2
rect 183 -3 184 -2
rect 184 -3 185 -2
rect 185 -3 186 -2
rect 186 -3 187 -2
rect 187 -3 188 -2
rect 188 -3 189 -2
rect 189 -3 190 -2
rect 190 -3 191 -2
rect 191 -3 192 -2
rect 192 -3 193 -2
rect 193 -3 194 -2
rect 194 -3 195 -2
rect 195 -3 196 -2
rect 196 -3 197 -2
rect 197 -3 198 -2
rect 198 -3 199 -2
rect 199 -3 200 -2
rect 200 -3 201 -2
rect 201 -3 202 -2
rect 202 -3 203 -2
rect 203 -3 204 -2
rect 204 -3 205 -2
rect 205 -3 206 -2
rect 206 -3 207 -2
rect 207 -3 208 -2
rect 208 -3 209 -2
rect 209 -3 210 -2
rect 210 -3 211 -2
rect 211 -3 212 -2
rect 212 -3 213 -2
rect 213 -3 214 -2
rect 214 -3 215 -2
rect 215 -3 216 -2
rect 216 -3 217 -2
rect 217 -3 218 -2
rect 218 -3 219 -2
rect 219 -3 220 -2
rect 220 -3 221 -2
rect 221 -3 222 -2
rect 222 -3 223 -2
rect 223 -3 224 -2
rect 224 -3 225 -2
rect 225 -3 226 -2
rect 226 -3 227 -2
rect 227 -3 228 -2
rect 228 -3 229 -2
rect 229 -3 230 -2
rect 230 -3 231 -2
rect 231 -3 232 -2
rect 232 -3 233 -2
rect 233 -3 234 -2
rect 234 -3 235 -2
rect 235 -3 236 -2
rect 236 -3 237 -2
rect 237 -3 238 -2
rect 238 -3 239 -2
rect 239 -3 240 -2
rect 240 -3 241 -2
rect 241 -3 242 -2
rect 242 -3 243 -2
rect 243 -3 244 -2
rect 244 -3 245 -2
rect 245 -3 246 -2
rect 246 -3 247 -2
rect 247 -3 248 -2
rect 248 -3 249 -2
rect 249 -3 250 -2
rect 250 -3 251 -2
rect 251 -3 252 -2
rect 252 -3 253 -2
rect 253 -3 254 -2
rect 254 -3 255 -2
rect 255 -3 256 -2
rect 256 -3 257 -2
rect 257 -3 258 -2
rect 258 -3 259 -2
rect 259 -3 260 -2
rect 260 -3 261 -2
rect 261 -3 262 -2
rect 262 -3 263 -2
rect 263 -3 264 -2
rect 264 -3 265 -2
rect 265 -3 266 -2
rect 266 -3 267 -2
rect 267 -3 268 -2
rect 268 -3 269 -2
rect 269 -3 270 -2
rect 270 -3 271 -2
rect 271 -3 272 -2
rect 272 -3 273 -2
rect 273 -3 274 -2
rect 274 -3 275 -2
rect 275 -3 276 -2
rect 276 -3 277 -2
rect 277 -3 278 -2
rect 278 -3 279 -2
rect 279 -3 280 -2
rect 280 -3 281 -2
rect 281 -3 282 -2
rect 282 -3 283 -2
rect 283 -3 284 -2
rect 284 -3 285 -2
rect 285 -3 286 -2
rect 286 -3 287 -2
rect 287 -3 288 -2
rect 288 -3 289 -2
rect 289 -3 290 -2
rect 290 -3 291 -2
rect 291 -3 292 -2
rect 292 -3 293 -2
rect 293 -3 294 -2
rect 294 -3 295 -2
rect 295 -3 296 -2
rect 296 -3 297 -2
rect 297 -3 298 -2
rect 298 -3 299 -2
rect 299 -3 300 -2
rect 300 -3 301 -2
rect 301 -3 302 -2
rect 302 -3 303 -2
rect 303 -3 304 -2
rect 304 -3 305 -2
rect 305 -3 306 -2
rect 306 -3 307 -2
rect 307 -3 308 -2
rect 308 -3 309 -2
rect 309 -3 310 -2
rect 310 -3 311 -2
rect 311 -3 312 -2
rect 312 -3 313 -2
rect 313 -3 314 -2
rect 314 -3 315 -2
rect 315 -3 316 -2
rect 316 -3 317 -2
rect 317 -3 318 -2
rect 318 -3 319 -2
rect 319 -3 320 -2
rect 320 -3 321 -2
rect 321 -3 322 -2
rect 322 -3 323 -2
rect 323 -3 324 -2
rect 324 -3 325 -2
rect 325 -3 326 -2
rect 326 -3 327 -2
rect 327 -3 328 -2
rect 328 -3 329 -2
rect 329 -3 330 -2
rect 330 -3 331 -2
rect 331 -3 332 -2
rect 332 -3 333 -2
rect 333 -3 334 -2
rect 334 -3 335 -2
rect 335 -3 336 -2
rect 336 -3 337 -2
rect 337 -3 338 -2
rect 338 -3 339 -2
rect 339 -3 340 -2
rect 340 -3 341 -2
rect 341 -3 342 -2
rect 342 -3 343 -2
rect 343 -3 344 -2
rect 344 -3 345 -2
rect 345 -3 346 -2
rect 346 -3 347 -2
rect 347 -3 348 -2
rect 348 -3 349 -2
rect 349 -3 350 -2
rect 350 -3 351 -2
rect 351 -3 352 -2
rect 352 -3 353 -2
rect 353 -3 354 -2
rect 354 -3 355 -2
rect 355 -3 356 -2
rect 356 -3 357 -2
rect 357 -3 358 -2
rect 358 -3 359 -2
rect 359 -3 360 -2
rect 360 -3 361 -2
rect 361 -3 362 -2
rect 362 -3 363 -2
rect 363 -3 364 -2
rect 364 -3 365 -2
rect 365 -3 366 -2
rect 366 -3 367 -2
rect 367 -3 368 -2
rect 368 -3 369 -2
rect 369 -3 370 -2
rect 370 -3 371 -2
rect 371 -3 372 -2
rect 372 -3 373 -2
rect 373 -3 374 -2
rect 374 -3 375 -2
rect 375 -3 376 -2
rect 376 -3 377 -2
rect 377 -3 378 -2
rect 378 -3 379 -2
rect 379 -3 380 -2
rect 380 -3 381 -2
rect 381 -3 382 -2
rect 382 -3 383 -2
rect 383 -3 384 -2
rect 384 -3 385 -2
rect 385 -3 386 -2
rect 386 -3 387 -2
rect 387 -3 388 -2
rect 388 -3 389 -2
rect 389 -3 390 -2
rect 390 -3 391 -2
rect 391 -3 392 -2
rect 392 -3 393 -2
rect 393 -3 394 -2
rect 394 -3 395 -2
rect 395 -3 396 -2
rect 396 -3 397 -2
rect 397 -3 398 -2
rect 398 -3 399 -2
rect 399 -3 400 -2
rect 400 -3 401 -2
rect 401 -3 402 -2
rect 402 -3 403 -2
rect 403 -3 404 -2
rect 404 -3 405 -2
rect 405 -3 406 -2
rect 406 -3 407 -2
rect 407 -3 408 -2
rect 408 -3 409 -2
rect 409 -3 410 -2
rect 410 -3 411 -2
rect 411 -3 412 -2
rect 412 -3 413 -2
rect 413 -3 414 -2
rect 414 -3 415 -2
rect 415 -3 416 -2
rect 416 -3 417 -2
rect 417 -3 418 -2
rect 418 -3 419 -2
rect 419 -3 420 -2
rect 420 -3 421 -2
rect 421 -3 422 -2
rect 422 -3 423 -2
rect 423 -3 424 -2
rect 424 -3 425 -2
rect 425 -3 426 -2
rect 426 -3 427 -2
rect 427 -3 428 -2
rect 428 -3 429 -2
rect 429 -3 430 -2
rect 430 -3 431 -2
rect 431 -3 432 -2
rect 432 -3 433 -2
rect 433 -3 434 -2
rect 434 -3 435 -2
rect 435 -3 436 -2
rect 436 -3 437 -2
rect 437 -3 438 -2
rect 438 -3 439 -2
rect 439 -3 440 -2
rect 440 -3 441 -2
rect 441 -3 442 -2
rect 442 -3 443 -2
rect 443 -3 444 -2
rect 444 -3 445 -2
rect 445 -3 446 -2
rect 446 -3 447 -2
rect 447 -3 448 -2
rect 448 -3 449 -2
rect 449 -3 450 -2
rect 450 -3 451 -2
rect 451 -3 452 -2
rect 452 -3 453 -2
rect 453 -3 454 -2
rect 454 -3 455 -2
rect 455 -3 456 -2
rect 456 -3 457 -2
rect 457 -3 458 -2
rect 458 -3 459 -2
rect 459 -3 460 -2
rect 460 -3 461 -2
rect 461 -3 462 -2
rect 462 -3 463 -2
rect 463 -3 464 -2
rect 464 -3 465 -2
rect 465 -3 466 -2
rect 466 -3 467 -2
rect 467 -3 468 -2
rect 468 -3 469 -2
rect 469 -3 470 -2
rect 470 -3 471 -2
rect 471 -3 472 -2
rect 472 -3 473 -2
rect 473 -3 474 -2
rect 474 -3 475 -2
rect 475 -3 476 -2
rect 476 -3 477 -2
rect 477 -3 478 -2
rect 478 -3 479 -2
rect 479 -3 480 -2
rect 2 -4 3 -3
rect 3 -4 4 -3
rect 4 -4 5 -3
rect 5 -4 6 -3
rect 6 -4 7 -3
rect 7 -4 8 -3
rect 8 -4 9 -3
rect 9 -4 10 -3
rect 10 -4 11 -3
rect 11 -4 12 -3
rect 12 -4 13 -3
rect 13 -4 14 -3
rect 14 -4 15 -3
rect 15 -4 16 -3
rect 16 -4 17 -3
rect 17 -4 18 -3
rect 18 -4 19 -3
rect 19 -4 20 -3
rect 20 -4 21 -3
rect 21 -4 22 -3
rect 22 -4 23 -3
rect 23 -4 24 -3
rect 24 -4 25 -3
rect 25 -4 26 -3
rect 26 -4 27 -3
rect 27 -4 28 -3
rect 28 -4 29 -3
rect 29 -4 30 -3
rect 30 -4 31 -3
rect 31 -4 32 -3
rect 32 -4 33 -3
rect 33 -4 34 -3
rect 34 -4 35 -3
rect 35 -4 36 -3
rect 36 -4 37 -3
rect 37 -4 38 -3
rect 38 -4 39 -3
rect 39 -4 40 -3
rect 40 -4 41 -3
rect 41 -4 42 -3
rect 42 -4 43 -3
rect 43 -4 44 -3
rect 44 -4 45 -3
rect 45 -4 46 -3
rect 46 -4 47 -3
rect 47 -4 48 -3
rect 48 -4 49 -3
rect 49 -4 50 -3
rect 50 -4 51 -3
rect 51 -4 52 -3
rect 52 -4 53 -3
rect 53 -4 54 -3
rect 54 -4 55 -3
rect 55 -4 56 -3
rect 56 -4 57 -3
rect 57 -4 58 -3
rect 58 -4 59 -3
rect 59 -4 60 -3
rect 60 -4 61 -3
rect 61 -4 62 -3
rect 62 -4 63 -3
rect 63 -4 64 -3
rect 64 -4 65 -3
rect 65 -4 66 -3
rect 66 -4 67 -3
rect 67 -4 68 -3
rect 68 -4 69 -3
rect 69 -4 70 -3
rect 70 -4 71 -3
rect 71 -4 72 -3
rect 72 -4 73 -3
rect 73 -4 74 -3
rect 74 -4 75 -3
rect 75 -4 76 -3
rect 76 -4 77 -3
rect 77 -4 78 -3
rect 78 -4 79 -3
rect 79 -4 80 -3
rect 80 -4 81 -3
rect 81 -4 82 -3
rect 82 -4 83 -3
rect 83 -4 84 -3
rect 84 -4 85 -3
rect 85 -4 86 -3
rect 86 -4 87 -3
rect 87 -4 88 -3
rect 88 -4 89 -3
rect 89 -4 90 -3
rect 90 -4 91 -3
rect 91 -4 92 -3
rect 92 -4 93 -3
rect 93 -4 94 -3
rect 94 -4 95 -3
rect 95 -4 96 -3
rect 96 -4 97 -3
rect 97 -4 98 -3
rect 98 -4 99 -3
rect 99 -4 100 -3
rect 100 -4 101 -3
rect 101 -4 102 -3
rect 102 -4 103 -3
rect 103 -4 104 -3
rect 104 -4 105 -3
rect 105 -4 106 -3
rect 106 -4 107 -3
rect 107 -4 108 -3
rect 108 -4 109 -3
rect 109 -4 110 -3
rect 110 -4 111 -3
rect 111 -4 112 -3
rect 112 -4 113 -3
rect 113 -4 114 -3
rect 114 -4 115 -3
rect 115 -4 116 -3
rect 116 -4 117 -3
rect 117 -4 118 -3
rect 118 -4 119 -3
rect 119 -4 120 -3
rect 120 -4 121 -3
rect 121 -4 122 -3
rect 122 -4 123 -3
rect 123 -4 124 -3
rect 124 -4 125 -3
rect 125 -4 126 -3
rect 126 -4 127 -3
rect 127 -4 128 -3
rect 128 -4 129 -3
rect 129 -4 130 -3
rect 130 -4 131 -3
rect 131 -4 132 -3
rect 132 -4 133 -3
rect 133 -4 134 -3
rect 134 -4 135 -3
rect 135 -4 136 -3
rect 136 -4 137 -3
rect 137 -4 138 -3
rect 138 -4 139 -3
rect 139 -4 140 -3
rect 140 -4 141 -3
rect 141 -4 142 -3
rect 142 -4 143 -3
rect 143 -4 144 -3
rect 144 -4 145 -3
rect 145 -4 146 -3
rect 146 -4 147 -3
rect 147 -4 148 -3
rect 148 -4 149 -3
rect 149 -4 150 -3
rect 150 -4 151 -3
rect 151 -4 152 -3
rect 152 -4 153 -3
rect 153 -4 154 -3
rect 154 -4 155 -3
rect 155 -4 156 -3
rect 156 -4 157 -3
rect 157 -4 158 -3
rect 158 -4 159 -3
rect 159 -4 160 -3
rect 160 -4 161 -3
rect 161 -4 162 -3
rect 162 -4 163 -3
rect 163 -4 164 -3
rect 164 -4 165 -3
rect 165 -4 166 -3
rect 166 -4 167 -3
rect 167 -4 168 -3
rect 168 -4 169 -3
rect 169 -4 170 -3
rect 170 -4 171 -3
rect 171 -4 172 -3
rect 172 -4 173 -3
rect 173 -4 174 -3
rect 174 -4 175 -3
rect 175 -4 176 -3
rect 176 -4 177 -3
rect 177 -4 178 -3
rect 178 -4 179 -3
rect 179 -4 180 -3
rect 180 -4 181 -3
rect 181 -4 182 -3
rect 182 -4 183 -3
rect 183 -4 184 -3
rect 184 -4 185 -3
rect 185 -4 186 -3
rect 186 -4 187 -3
rect 187 -4 188 -3
rect 188 -4 189 -3
rect 189 -4 190 -3
rect 190 -4 191 -3
rect 191 -4 192 -3
rect 192 -4 193 -3
rect 193 -4 194 -3
rect 194 -4 195 -3
rect 195 -4 196 -3
rect 196 -4 197 -3
rect 197 -4 198 -3
rect 198 -4 199 -3
rect 199 -4 200 -3
rect 200 -4 201 -3
rect 201 -4 202 -3
rect 202 -4 203 -3
rect 203 -4 204 -3
rect 204 -4 205 -3
rect 205 -4 206 -3
rect 206 -4 207 -3
rect 207 -4 208 -3
rect 208 -4 209 -3
rect 209 -4 210 -3
rect 210 -4 211 -3
rect 211 -4 212 -3
rect 212 -4 213 -3
rect 213 -4 214 -3
rect 214 -4 215 -3
rect 215 -4 216 -3
rect 216 -4 217 -3
rect 217 -4 218 -3
rect 218 -4 219 -3
rect 219 -4 220 -3
rect 220 -4 221 -3
rect 221 -4 222 -3
rect 222 -4 223 -3
rect 223 -4 224 -3
rect 224 -4 225 -3
rect 225 -4 226 -3
rect 226 -4 227 -3
rect 227 -4 228 -3
rect 228 -4 229 -3
rect 229 -4 230 -3
rect 230 -4 231 -3
rect 231 -4 232 -3
rect 232 -4 233 -3
rect 233 -4 234 -3
rect 234 -4 235 -3
rect 235 -4 236 -3
rect 236 -4 237 -3
rect 237 -4 238 -3
rect 238 -4 239 -3
rect 239 -4 240 -3
rect 240 -4 241 -3
rect 241 -4 242 -3
rect 242 -4 243 -3
rect 243 -4 244 -3
rect 244 -4 245 -3
rect 245 -4 246 -3
rect 246 -4 247 -3
rect 247 -4 248 -3
rect 248 -4 249 -3
rect 249 -4 250 -3
rect 250 -4 251 -3
rect 251 -4 252 -3
rect 252 -4 253 -3
rect 253 -4 254 -3
rect 254 -4 255 -3
rect 255 -4 256 -3
rect 256 -4 257 -3
rect 257 -4 258 -3
rect 258 -4 259 -3
rect 259 -4 260 -3
rect 260 -4 261 -3
rect 261 -4 262 -3
rect 262 -4 263 -3
rect 263 -4 264 -3
rect 264 -4 265 -3
rect 265 -4 266 -3
rect 266 -4 267 -3
rect 267 -4 268 -3
rect 268 -4 269 -3
rect 269 -4 270 -3
rect 270 -4 271 -3
rect 271 -4 272 -3
rect 272 -4 273 -3
rect 273 -4 274 -3
rect 274 -4 275 -3
rect 275 -4 276 -3
rect 276 -4 277 -3
rect 277 -4 278 -3
rect 278 -4 279 -3
rect 279 -4 280 -3
rect 280 -4 281 -3
rect 281 -4 282 -3
rect 282 -4 283 -3
rect 283 -4 284 -3
rect 284 -4 285 -3
rect 285 -4 286 -3
rect 286 -4 287 -3
rect 287 -4 288 -3
rect 288 -4 289 -3
rect 289 -4 290 -3
rect 290 -4 291 -3
rect 291 -4 292 -3
rect 292 -4 293 -3
rect 293 -4 294 -3
rect 294 -4 295 -3
rect 295 -4 296 -3
rect 296 -4 297 -3
rect 297 -4 298 -3
rect 298 -4 299 -3
rect 299 -4 300 -3
rect 300 -4 301 -3
rect 301 -4 302 -3
rect 302 -4 303 -3
rect 303 -4 304 -3
rect 304 -4 305 -3
rect 305 -4 306 -3
rect 306 -4 307 -3
rect 307 -4 308 -3
rect 308 -4 309 -3
rect 309 -4 310 -3
rect 310 -4 311 -3
rect 311 -4 312 -3
rect 312 -4 313 -3
rect 313 -4 314 -3
rect 314 -4 315 -3
rect 315 -4 316 -3
rect 316 -4 317 -3
rect 317 -4 318 -3
rect 318 -4 319 -3
rect 319 -4 320 -3
rect 320 -4 321 -3
rect 321 -4 322 -3
rect 322 -4 323 -3
rect 323 -4 324 -3
rect 324 -4 325 -3
rect 325 -4 326 -3
rect 326 -4 327 -3
rect 327 -4 328 -3
rect 328 -4 329 -3
rect 329 -4 330 -3
rect 330 -4 331 -3
rect 331 -4 332 -3
rect 332 -4 333 -3
rect 333 -4 334 -3
rect 334 -4 335 -3
rect 335 -4 336 -3
rect 336 -4 337 -3
rect 337 -4 338 -3
rect 338 -4 339 -3
rect 339 -4 340 -3
rect 340 -4 341 -3
rect 341 -4 342 -3
rect 342 -4 343 -3
rect 343 -4 344 -3
rect 344 -4 345 -3
rect 345 -4 346 -3
rect 346 -4 347 -3
rect 347 -4 348 -3
rect 348 -4 349 -3
rect 349 -4 350 -3
rect 350 -4 351 -3
rect 351 -4 352 -3
rect 352 -4 353 -3
rect 353 -4 354 -3
rect 354 -4 355 -3
rect 355 -4 356 -3
rect 356 -4 357 -3
rect 357 -4 358 -3
rect 358 -4 359 -3
rect 359 -4 360 -3
rect 360 -4 361 -3
rect 361 -4 362 -3
rect 362 -4 363 -3
rect 363 -4 364 -3
rect 364 -4 365 -3
rect 365 -4 366 -3
rect 366 -4 367 -3
rect 367 -4 368 -3
rect 368 -4 369 -3
rect 369 -4 370 -3
rect 370 -4 371 -3
rect 371 -4 372 -3
rect 372 -4 373 -3
rect 373 -4 374 -3
rect 374 -4 375 -3
rect 375 -4 376 -3
rect 376 -4 377 -3
rect 377 -4 378 -3
rect 378 -4 379 -3
rect 379 -4 380 -3
rect 380 -4 381 -3
rect 381 -4 382 -3
rect 382 -4 383 -3
rect 383 -4 384 -3
rect 384 -4 385 -3
rect 385 -4 386 -3
rect 386 -4 387 -3
rect 387 -4 388 -3
rect 388 -4 389 -3
rect 389 -4 390 -3
rect 390 -4 391 -3
rect 391 -4 392 -3
rect 392 -4 393 -3
rect 393 -4 394 -3
rect 394 -4 395 -3
rect 395 -4 396 -3
rect 396 -4 397 -3
rect 397 -4 398 -3
rect 398 -4 399 -3
rect 399 -4 400 -3
rect 400 -4 401 -3
rect 401 -4 402 -3
rect 402 -4 403 -3
rect 403 -4 404 -3
rect 404 -4 405 -3
rect 405 -4 406 -3
rect 406 -4 407 -3
rect 407 -4 408 -3
rect 408 -4 409 -3
rect 409 -4 410 -3
rect 410 -4 411 -3
rect 411 -4 412 -3
rect 412 -4 413 -3
rect 413 -4 414 -3
rect 414 -4 415 -3
rect 415 -4 416 -3
rect 416 -4 417 -3
rect 417 -4 418 -3
rect 418 -4 419 -3
rect 419 -4 420 -3
rect 420 -4 421 -3
rect 421 -4 422 -3
rect 422 -4 423 -3
rect 423 -4 424 -3
rect 424 -4 425 -3
rect 425 -4 426 -3
rect 426 -4 427 -3
rect 427 -4 428 -3
rect 428 -4 429 -3
rect 429 -4 430 -3
rect 430 -4 431 -3
rect 431 -4 432 -3
rect 432 -4 433 -3
rect 433 -4 434 -3
rect 434 -4 435 -3
rect 435 -4 436 -3
rect 436 -4 437 -3
rect 437 -4 438 -3
rect 438 -4 439 -3
rect 439 -4 440 -3
rect 440 -4 441 -3
rect 441 -4 442 -3
rect 442 -4 443 -3
rect 443 -4 444 -3
rect 444 -4 445 -3
rect 445 -4 446 -3
rect 446 -4 447 -3
rect 447 -4 448 -3
rect 448 -4 449 -3
rect 449 -4 450 -3
rect 450 -4 451 -3
rect 451 -4 452 -3
rect 452 -4 453 -3
rect 453 -4 454 -3
rect 454 -4 455 -3
rect 455 -4 456 -3
rect 456 -4 457 -3
rect 457 -4 458 -3
rect 458 -4 459 -3
rect 459 -4 460 -3
rect 460 -4 461 -3
rect 461 -4 462 -3
rect 462 -4 463 -3
rect 463 -4 464 -3
rect 464 -4 465 -3
rect 465 -4 466 -3
rect 466 -4 467 -3
rect 467 -4 468 -3
rect 468 -4 469 -3
rect 469 -4 470 -3
rect 470 -4 471 -3
rect 471 -4 472 -3
rect 472 -4 473 -3
rect 473 -4 474 -3
rect 474 -4 475 -3
rect 475 -4 476 -3
rect 476 -4 477 -3
rect 477 -4 478 -3
rect 478 -4 479 -3
rect 479 -4 480 -3
rect 2 -5 3 -4
rect 3 -5 4 -4
rect 4 -5 5 -4
rect 5 -5 6 -4
rect 6 -5 7 -4
rect 7 -5 8 -4
rect 8 -5 9 -4
rect 9 -5 10 -4
rect 10 -5 11 -4
rect 11 -5 12 -4
rect 12 -5 13 -4
rect 13 -5 14 -4
rect 14 -5 15 -4
rect 15 -5 16 -4
rect 16 -5 17 -4
rect 17 -5 18 -4
rect 18 -5 19 -4
rect 19 -5 20 -4
rect 20 -5 21 -4
rect 21 -5 22 -4
rect 22 -5 23 -4
rect 23 -5 24 -4
rect 24 -5 25 -4
rect 25 -5 26 -4
rect 26 -5 27 -4
rect 27 -5 28 -4
rect 28 -5 29 -4
rect 29 -5 30 -4
rect 30 -5 31 -4
rect 31 -5 32 -4
rect 32 -5 33 -4
rect 33 -5 34 -4
rect 34 -5 35 -4
rect 35 -5 36 -4
rect 36 -5 37 -4
rect 37 -5 38 -4
rect 38 -5 39 -4
rect 39 -5 40 -4
rect 40 -5 41 -4
rect 41 -5 42 -4
rect 42 -5 43 -4
rect 43 -5 44 -4
rect 44 -5 45 -4
rect 45 -5 46 -4
rect 46 -5 47 -4
rect 47 -5 48 -4
rect 48 -5 49 -4
rect 49 -5 50 -4
rect 50 -5 51 -4
rect 51 -5 52 -4
rect 52 -5 53 -4
rect 53 -5 54 -4
rect 54 -5 55 -4
rect 55 -5 56 -4
rect 56 -5 57 -4
rect 57 -5 58 -4
rect 58 -5 59 -4
rect 59 -5 60 -4
rect 60 -5 61 -4
rect 61 -5 62 -4
rect 62 -5 63 -4
rect 63 -5 64 -4
rect 64 -5 65 -4
rect 65 -5 66 -4
rect 66 -5 67 -4
rect 67 -5 68 -4
rect 68 -5 69 -4
rect 69 -5 70 -4
rect 70 -5 71 -4
rect 71 -5 72 -4
rect 72 -5 73 -4
rect 73 -5 74 -4
rect 74 -5 75 -4
rect 75 -5 76 -4
rect 76 -5 77 -4
rect 77 -5 78 -4
rect 78 -5 79 -4
rect 79 -5 80 -4
rect 80 -5 81 -4
rect 81 -5 82 -4
rect 82 -5 83 -4
rect 83 -5 84 -4
rect 84 -5 85 -4
rect 85 -5 86 -4
rect 86 -5 87 -4
rect 87 -5 88 -4
rect 88 -5 89 -4
rect 89 -5 90 -4
rect 90 -5 91 -4
rect 91 -5 92 -4
rect 92 -5 93 -4
rect 93 -5 94 -4
rect 94 -5 95 -4
rect 95 -5 96 -4
rect 96 -5 97 -4
rect 97 -5 98 -4
rect 98 -5 99 -4
rect 99 -5 100 -4
rect 100 -5 101 -4
rect 101 -5 102 -4
rect 102 -5 103 -4
rect 103 -5 104 -4
rect 104 -5 105 -4
rect 105 -5 106 -4
rect 106 -5 107 -4
rect 107 -5 108 -4
rect 108 -5 109 -4
rect 109 -5 110 -4
rect 110 -5 111 -4
rect 111 -5 112 -4
rect 112 -5 113 -4
rect 113 -5 114 -4
rect 114 -5 115 -4
rect 115 -5 116 -4
rect 116 -5 117 -4
rect 117 -5 118 -4
rect 118 -5 119 -4
rect 119 -5 120 -4
rect 120 -5 121 -4
rect 121 -5 122 -4
rect 122 -5 123 -4
rect 123 -5 124 -4
rect 124 -5 125 -4
rect 125 -5 126 -4
rect 126 -5 127 -4
rect 127 -5 128 -4
rect 128 -5 129 -4
rect 129 -5 130 -4
rect 130 -5 131 -4
rect 131 -5 132 -4
rect 132 -5 133 -4
rect 133 -5 134 -4
rect 134 -5 135 -4
rect 135 -5 136 -4
rect 136 -5 137 -4
rect 137 -5 138 -4
rect 138 -5 139 -4
rect 139 -5 140 -4
rect 140 -5 141 -4
rect 141 -5 142 -4
rect 142 -5 143 -4
rect 143 -5 144 -4
rect 144 -5 145 -4
rect 145 -5 146 -4
rect 146 -5 147 -4
rect 147 -5 148 -4
rect 148 -5 149 -4
rect 149 -5 150 -4
rect 150 -5 151 -4
rect 151 -5 152 -4
rect 152 -5 153 -4
rect 153 -5 154 -4
rect 154 -5 155 -4
rect 155 -5 156 -4
rect 156 -5 157 -4
rect 157 -5 158 -4
rect 158 -5 159 -4
rect 159 -5 160 -4
rect 160 -5 161 -4
rect 161 -5 162 -4
rect 162 -5 163 -4
rect 163 -5 164 -4
rect 164 -5 165 -4
rect 165 -5 166 -4
rect 166 -5 167 -4
rect 167 -5 168 -4
rect 168 -5 169 -4
rect 169 -5 170 -4
rect 170 -5 171 -4
rect 171 -5 172 -4
rect 172 -5 173 -4
rect 173 -5 174 -4
rect 174 -5 175 -4
rect 175 -5 176 -4
rect 176 -5 177 -4
rect 177 -5 178 -4
rect 178 -5 179 -4
rect 179 -5 180 -4
rect 180 -5 181 -4
rect 181 -5 182 -4
rect 182 -5 183 -4
rect 183 -5 184 -4
rect 184 -5 185 -4
rect 185 -5 186 -4
rect 186 -5 187 -4
rect 187 -5 188 -4
rect 188 -5 189 -4
rect 189 -5 190 -4
rect 190 -5 191 -4
rect 191 -5 192 -4
rect 192 -5 193 -4
rect 193 -5 194 -4
rect 194 -5 195 -4
rect 195 -5 196 -4
rect 196 -5 197 -4
rect 197 -5 198 -4
rect 198 -5 199 -4
rect 199 -5 200 -4
rect 200 -5 201 -4
rect 201 -5 202 -4
rect 202 -5 203 -4
rect 203 -5 204 -4
rect 204 -5 205 -4
rect 205 -5 206 -4
rect 206 -5 207 -4
rect 207 -5 208 -4
rect 208 -5 209 -4
rect 209 -5 210 -4
rect 210 -5 211 -4
rect 211 -5 212 -4
rect 212 -5 213 -4
rect 213 -5 214 -4
rect 214 -5 215 -4
rect 215 -5 216 -4
rect 216 -5 217 -4
rect 217 -5 218 -4
rect 218 -5 219 -4
rect 219 -5 220 -4
rect 220 -5 221 -4
rect 221 -5 222 -4
rect 222 -5 223 -4
rect 223 -5 224 -4
rect 224 -5 225 -4
rect 225 -5 226 -4
rect 226 -5 227 -4
rect 227 -5 228 -4
rect 228 -5 229 -4
rect 229 -5 230 -4
rect 230 -5 231 -4
rect 231 -5 232 -4
rect 232 -5 233 -4
rect 233 -5 234 -4
rect 234 -5 235 -4
rect 235 -5 236 -4
rect 236 -5 237 -4
rect 237 -5 238 -4
rect 238 -5 239 -4
rect 239 -5 240 -4
rect 240 -5 241 -4
rect 241 -5 242 -4
rect 242 -5 243 -4
rect 243 -5 244 -4
rect 244 -5 245 -4
rect 245 -5 246 -4
rect 246 -5 247 -4
rect 247 -5 248 -4
rect 248 -5 249 -4
rect 249 -5 250 -4
rect 250 -5 251 -4
rect 251 -5 252 -4
rect 252 -5 253 -4
rect 253 -5 254 -4
rect 254 -5 255 -4
rect 255 -5 256 -4
rect 256 -5 257 -4
rect 257 -5 258 -4
rect 258 -5 259 -4
rect 259 -5 260 -4
rect 260 -5 261 -4
rect 261 -5 262 -4
rect 262 -5 263 -4
rect 263 -5 264 -4
rect 264 -5 265 -4
rect 265 -5 266 -4
rect 266 -5 267 -4
rect 267 -5 268 -4
rect 268 -5 269 -4
rect 269 -5 270 -4
rect 270 -5 271 -4
rect 271 -5 272 -4
rect 272 -5 273 -4
rect 273 -5 274 -4
rect 274 -5 275 -4
rect 275 -5 276 -4
rect 276 -5 277 -4
rect 277 -5 278 -4
rect 278 -5 279 -4
rect 279 -5 280 -4
rect 280 -5 281 -4
rect 281 -5 282 -4
rect 282 -5 283 -4
rect 283 -5 284 -4
rect 284 -5 285 -4
rect 285 -5 286 -4
rect 286 -5 287 -4
rect 287 -5 288 -4
rect 288 -5 289 -4
rect 289 -5 290 -4
rect 290 -5 291 -4
rect 291 -5 292 -4
rect 292 -5 293 -4
rect 293 -5 294 -4
rect 294 -5 295 -4
rect 295 -5 296 -4
rect 296 -5 297 -4
rect 297 -5 298 -4
rect 298 -5 299 -4
rect 299 -5 300 -4
rect 300 -5 301 -4
rect 301 -5 302 -4
rect 302 -5 303 -4
rect 303 -5 304 -4
rect 304 -5 305 -4
rect 305 -5 306 -4
rect 306 -5 307 -4
rect 307 -5 308 -4
rect 308 -5 309 -4
rect 309 -5 310 -4
rect 310 -5 311 -4
rect 311 -5 312 -4
rect 312 -5 313 -4
rect 313 -5 314 -4
rect 314 -5 315 -4
rect 315 -5 316 -4
rect 316 -5 317 -4
rect 317 -5 318 -4
rect 318 -5 319 -4
rect 319 -5 320 -4
rect 320 -5 321 -4
rect 321 -5 322 -4
rect 322 -5 323 -4
rect 323 -5 324 -4
rect 324 -5 325 -4
rect 325 -5 326 -4
rect 326 -5 327 -4
rect 327 -5 328 -4
rect 328 -5 329 -4
rect 329 -5 330 -4
rect 330 -5 331 -4
rect 331 -5 332 -4
rect 332 -5 333 -4
rect 333 -5 334 -4
rect 334 -5 335 -4
rect 335 -5 336 -4
rect 336 -5 337 -4
rect 337 -5 338 -4
rect 338 -5 339 -4
rect 339 -5 340 -4
rect 340 -5 341 -4
rect 341 -5 342 -4
rect 342 -5 343 -4
rect 343 -5 344 -4
rect 344 -5 345 -4
rect 345 -5 346 -4
rect 346 -5 347 -4
rect 347 -5 348 -4
rect 348 -5 349 -4
rect 349 -5 350 -4
rect 350 -5 351 -4
rect 351 -5 352 -4
rect 352 -5 353 -4
rect 353 -5 354 -4
rect 354 -5 355 -4
rect 355 -5 356 -4
rect 356 -5 357 -4
rect 357 -5 358 -4
rect 358 -5 359 -4
rect 359 -5 360 -4
rect 360 -5 361 -4
rect 361 -5 362 -4
rect 362 -5 363 -4
rect 363 -5 364 -4
rect 364 -5 365 -4
rect 365 -5 366 -4
rect 366 -5 367 -4
rect 367 -5 368 -4
rect 368 -5 369 -4
rect 369 -5 370 -4
rect 370 -5 371 -4
rect 371 -5 372 -4
rect 372 -5 373 -4
rect 373 -5 374 -4
rect 374 -5 375 -4
rect 375 -5 376 -4
rect 376 -5 377 -4
rect 377 -5 378 -4
rect 378 -5 379 -4
rect 379 -5 380 -4
rect 380 -5 381 -4
rect 381 -5 382 -4
rect 382 -5 383 -4
rect 383 -5 384 -4
rect 384 -5 385 -4
rect 385 -5 386 -4
rect 386 -5 387 -4
rect 387 -5 388 -4
rect 388 -5 389 -4
rect 389 -5 390 -4
rect 390 -5 391 -4
rect 391 -5 392 -4
rect 392 -5 393 -4
rect 393 -5 394 -4
rect 394 -5 395 -4
rect 395 -5 396 -4
rect 396 -5 397 -4
rect 397 -5 398 -4
rect 398 -5 399 -4
rect 399 -5 400 -4
rect 400 -5 401 -4
rect 401 -5 402 -4
rect 402 -5 403 -4
rect 403 -5 404 -4
rect 404 -5 405 -4
rect 405 -5 406 -4
rect 406 -5 407 -4
rect 407 -5 408 -4
rect 408 -5 409 -4
rect 409 -5 410 -4
rect 410 -5 411 -4
rect 411 -5 412 -4
rect 412 -5 413 -4
rect 413 -5 414 -4
rect 414 -5 415 -4
rect 415 -5 416 -4
rect 416 -5 417 -4
rect 417 -5 418 -4
rect 418 -5 419 -4
rect 419 -5 420 -4
rect 420 -5 421 -4
rect 421 -5 422 -4
rect 422 -5 423 -4
rect 423 -5 424 -4
rect 424 -5 425 -4
rect 425 -5 426 -4
rect 426 -5 427 -4
rect 427 -5 428 -4
rect 428 -5 429 -4
rect 429 -5 430 -4
rect 430 -5 431 -4
rect 431 -5 432 -4
rect 432 -5 433 -4
rect 433 -5 434 -4
rect 434 -5 435 -4
rect 435 -5 436 -4
rect 436 -5 437 -4
rect 437 -5 438 -4
rect 438 -5 439 -4
rect 439 -5 440 -4
rect 440 -5 441 -4
rect 441 -5 442 -4
rect 442 -5 443 -4
rect 443 -5 444 -4
rect 444 -5 445 -4
rect 445 -5 446 -4
rect 446 -5 447 -4
rect 447 -5 448 -4
rect 448 -5 449 -4
rect 449 -5 450 -4
rect 450 -5 451 -4
rect 451 -5 452 -4
rect 452 -5 453 -4
rect 453 -5 454 -4
rect 454 -5 455 -4
rect 455 -5 456 -4
rect 456 -5 457 -4
rect 457 -5 458 -4
rect 458 -5 459 -4
rect 459 -5 460 -4
rect 460 -5 461 -4
rect 461 -5 462 -4
rect 462 -5 463 -4
rect 463 -5 464 -4
rect 464 -5 465 -4
rect 465 -5 466 -4
rect 466 -5 467 -4
rect 467 -5 468 -4
rect 468 -5 469 -4
rect 469 -5 470 -4
rect 470 -5 471 -4
rect 471 -5 472 -4
rect 472 -5 473 -4
rect 473 -5 474 -4
rect 474 -5 475 -4
rect 475 -5 476 -4
rect 476 -5 477 -4
rect 477 -5 478 -4
rect 478 -5 479 -4
rect 479 -5 480 -4
rect 2 -6 3 -5
rect 3 -6 4 -5
rect 4 -6 5 -5
rect 5 -6 6 -5
rect 6 -6 7 -5
rect 7 -6 8 -5
rect 8 -6 9 -5
rect 9 -6 10 -5
rect 10 -6 11 -5
rect 11 -6 12 -5
rect 12 -6 13 -5
rect 13 -6 14 -5
rect 14 -6 15 -5
rect 18 -6 19 -5
rect 19 -6 20 -5
rect 20 -6 21 -5
rect 21 -6 22 -5
rect 22 -6 23 -5
rect 23 -6 24 -5
rect 24 -6 25 -5
rect 25 -6 26 -5
rect 26 -6 27 -5
rect 27 -6 28 -5
rect 28 -6 29 -5
rect 29 -6 30 -5
rect 30 -6 31 -5
rect 31 -6 32 -5
rect 32 -6 33 -5
rect 33 -6 34 -5
rect 34 -6 35 -5
rect 35 -6 36 -5
rect 36 -6 37 -5
rect 37 -6 38 -5
rect 38 -6 39 -5
rect 39 -6 40 -5
rect 40 -6 41 -5
rect 41 -6 42 -5
rect 42 -6 43 -5
rect 43 -6 44 -5
rect 44 -6 45 -5
rect 45 -6 46 -5
rect 46 -6 47 -5
rect 50 -6 51 -5
rect 51 -6 52 -5
rect 52 -6 53 -5
rect 53 -6 54 -5
rect 54 -6 55 -5
rect 55 -6 56 -5
rect 56 -6 57 -5
rect 57 -6 58 -5
rect 58 -6 59 -5
rect 59 -6 60 -5
rect 60 -6 61 -5
rect 61 -6 62 -5
rect 62 -6 63 -5
rect 63 -6 64 -5
rect 64 -6 65 -5
rect 65 -6 66 -5
rect 66 -6 67 -5
rect 67 -6 68 -5
rect 68 -6 69 -5
rect 69 -6 70 -5
rect 70 -6 71 -5
rect 71 -6 72 -5
rect 72 -6 73 -5
rect 73 -6 74 -5
rect 74 -6 75 -5
rect 75 -6 76 -5
rect 76 -6 77 -5
rect 77 -6 78 -5
rect 78 -6 79 -5
rect 82 -6 83 -5
rect 83 -6 84 -5
rect 84 -6 85 -5
rect 85 -6 86 -5
rect 86 -6 87 -5
rect 87 -6 88 -5
rect 88 -6 89 -5
rect 89 -6 90 -5
rect 90 -6 91 -5
rect 91 -6 92 -5
rect 92 -6 93 -5
rect 93 -6 94 -5
rect 94 -6 95 -5
rect 95 -6 96 -5
rect 96 -6 97 -5
rect 97 -6 98 -5
rect 98 -6 99 -5
rect 99 -6 100 -5
rect 100 -6 101 -5
rect 101 -6 102 -5
rect 102 -6 103 -5
rect 103 -6 104 -5
rect 104 -6 105 -5
rect 105 -6 106 -5
rect 106 -6 107 -5
rect 107 -6 108 -5
rect 108 -6 109 -5
rect 109 -6 110 -5
rect 110 -6 111 -5
rect 114 -6 115 -5
rect 115 -6 116 -5
rect 116 -6 117 -5
rect 117 -6 118 -5
rect 118 -6 119 -5
rect 119 -6 120 -5
rect 120 -6 121 -5
rect 121 -6 122 -5
rect 122 -6 123 -5
rect 123 -6 124 -5
rect 124 -6 125 -5
rect 125 -6 126 -5
rect 126 -6 127 -5
rect 127 -6 128 -5
rect 128 -6 129 -5
rect 129 -6 130 -5
rect 130 -6 131 -5
rect 131 -6 132 -5
rect 132 -6 133 -5
rect 133 -6 134 -5
rect 134 -6 135 -5
rect 135 -6 136 -5
rect 136 -6 137 -5
rect 137 -6 138 -5
rect 138 -6 139 -5
rect 139 -6 140 -5
rect 140 -6 141 -5
rect 141 -6 142 -5
rect 142 -6 143 -5
rect 146 -6 147 -5
rect 147 -6 148 -5
rect 148 -6 149 -5
rect 149 -6 150 -5
rect 150 -6 151 -5
rect 151 -6 152 -5
rect 152 -6 153 -5
rect 153 -6 154 -5
rect 154 -6 155 -5
rect 155 -6 156 -5
rect 156 -6 157 -5
rect 157 -6 158 -5
rect 158 -6 159 -5
rect 159 -6 160 -5
rect 160 -6 161 -5
rect 161 -6 162 -5
rect 162 -6 163 -5
rect 163 -6 164 -5
rect 164 -6 165 -5
rect 165 -6 166 -5
rect 166 -6 167 -5
rect 167 -6 168 -5
rect 168 -6 169 -5
rect 169 -6 170 -5
rect 170 -6 171 -5
rect 171 -6 172 -5
rect 172 -6 173 -5
rect 173 -6 174 -5
rect 174 -6 175 -5
rect 178 -6 179 -5
rect 179 -6 180 -5
rect 180 -6 181 -5
rect 181 -6 182 -5
rect 182 -6 183 -5
rect 183 -6 184 -5
rect 184 -6 185 -5
rect 185 -6 186 -5
rect 186 -6 187 -5
rect 187 -6 188 -5
rect 188 -6 189 -5
rect 189 -6 190 -5
rect 190 -6 191 -5
rect 191 -6 192 -5
rect 192 -6 193 -5
rect 193 -6 194 -5
rect 194 -6 195 -5
rect 195 -6 196 -5
rect 196 -6 197 -5
rect 197 -6 198 -5
rect 198 -6 199 -5
rect 199 -6 200 -5
rect 200 -6 201 -5
rect 201 -6 202 -5
rect 202 -6 203 -5
rect 203 -6 204 -5
rect 204 -6 205 -5
rect 205 -6 206 -5
rect 206 -6 207 -5
rect 207 -6 208 -5
rect 208 -6 209 -5
rect 209 -6 210 -5
rect 210 -6 211 -5
rect 211 -6 212 -5
rect 212 -6 213 -5
rect 213 -6 214 -5
rect 214 -6 215 -5
rect 215 -6 216 -5
rect 216 -6 217 -5
rect 217 -6 218 -5
rect 218 -6 219 -5
rect 219 -6 220 -5
rect 220 -6 221 -5
rect 221 -6 222 -5
rect 222 -6 223 -5
rect 223 -6 224 -5
rect 224 -6 225 -5
rect 225 -6 226 -5
rect 226 -6 227 -5
rect 227 -6 228 -5
rect 228 -6 229 -5
rect 229 -6 230 -5
rect 230 -6 231 -5
rect 231 -6 232 -5
rect 232 -6 233 -5
rect 233 -6 234 -5
rect 234 -6 235 -5
rect 235 -6 236 -5
rect 236 -6 237 -5
rect 237 -6 238 -5
rect 238 -6 239 -5
rect 239 -6 240 -5
rect 240 -6 241 -5
rect 241 -6 242 -5
rect 242 -6 243 -5
rect 243 -6 244 -5
rect 244 -6 245 -5
rect 245 -6 246 -5
rect 246 -6 247 -5
rect 247 -6 248 -5
rect 248 -6 249 -5
rect 249 -6 250 -5
rect 250 -6 251 -5
rect 251 -6 252 -5
rect 252 -6 253 -5
rect 253 -6 254 -5
rect 254 -6 255 -5
rect 255 -6 256 -5
rect 256 -6 257 -5
rect 257 -6 258 -5
rect 258 -6 259 -5
rect 259 -6 260 -5
rect 260 -6 261 -5
rect 261 -6 262 -5
rect 262 -6 263 -5
rect 263 -6 264 -5
rect 264 -6 265 -5
rect 265 -6 266 -5
rect 266 -6 267 -5
rect 267 -6 268 -5
rect 268 -6 269 -5
rect 269 -6 270 -5
rect 270 -6 271 -5
rect 271 -6 272 -5
rect 272 -6 273 -5
rect 273 -6 274 -5
rect 274 -6 275 -5
rect 275 -6 276 -5
rect 276 -6 277 -5
rect 277 -6 278 -5
rect 278 -6 279 -5
rect 279 -6 280 -5
rect 280 -6 281 -5
rect 281 -6 282 -5
rect 282 -6 283 -5
rect 283 -6 284 -5
rect 284 -6 285 -5
rect 285 -6 286 -5
rect 286 -6 287 -5
rect 287 -6 288 -5
rect 288 -6 289 -5
rect 289 -6 290 -5
rect 290 -6 291 -5
rect 291 -6 292 -5
rect 292 -6 293 -5
rect 293 -6 294 -5
rect 294 -6 295 -5
rect 295 -6 296 -5
rect 296 -6 297 -5
rect 297 -6 298 -5
rect 298 -6 299 -5
rect 299 -6 300 -5
rect 300 -6 301 -5
rect 301 -6 302 -5
rect 302 -6 303 -5
rect 303 -6 304 -5
rect 304 -6 305 -5
rect 305 -6 306 -5
rect 306 -6 307 -5
rect 307 -6 308 -5
rect 308 -6 309 -5
rect 309 -6 310 -5
rect 310 -6 311 -5
rect 311 -6 312 -5
rect 312 -6 313 -5
rect 313 -6 314 -5
rect 314 -6 315 -5
rect 315 -6 316 -5
rect 316 -6 317 -5
rect 317 -6 318 -5
rect 318 -6 319 -5
rect 319 -6 320 -5
rect 320 -6 321 -5
rect 321 -6 322 -5
rect 322 -6 323 -5
rect 323 -6 324 -5
rect 324 -6 325 -5
rect 325 -6 326 -5
rect 326 -6 327 -5
rect 327 -6 328 -5
rect 328 -6 329 -5
rect 329 -6 330 -5
rect 330 -6 331 -5
rect 331 -6 332 -5
rect 332 -6 333 -5
rect 333 -6 334 -5
rect 334 -6 335 -5
rect 335 -6 336 -5
rect 336 -6 337 -5
rect 337 -6 338 -5
rect 338 -6 339 -5
rect 339 -6 340 -5
rect 340 -6 341 -5
rect 341 -6 342 -5
rect 342 -6 343 -5
rect 343 -6 344 -5
rect 344 -6 345 -5
rect 345 -6 346 -5
rect 346 -6 347 -5
rect 347 -6 348 -5
rect 348 -6 349 -5
rect 349 -6 350 -5
rect 350 -6 351 -5
rect 351 -6 352 -5
rect 352 -6 353 -5
rect 353 -6 354 -5
rect 354 -6 355 -5
rect 355 -6 356 -5
rect 356 -6 357 -5
rect 357 -6 358 -5
rect 358 -6 359 -5
rect 359 -6 360 -5
rect 360 -6 361 -5
rect 361 -6 362 -5
rect 362 -6 363 -5
rect 363 -6 364 -5
rect 364 -6 365 -5
rect 365 -6 366 -5
rect 366 -6 367 -5
rect 367 -6 368 -5
rect 368 -6 369 -5
rect 369 -6 370 -5
rect 370 -6 371 -5
rect 371 -6 372 -5
rect 372 -6 373 -5
rect 373 -6 374 -5
rect 374 -6 375 -5
rect 375 -6 376 -5
rect 376 -6 377 -5
rect 377 -6 378 -5
rect 378 -6 379 -5
rect 379 -6 380 -5
rect 380 -6 381 -5
rect 381 -6 382 -5
rect 382 -6 383 -5
rect 383 -6 384 -5
rect 384 -6 385 -5
rect 385 -6 386 -5
rect 386 -6 387 -5
rect 387 -6 388 -5
rect 388 -6 389 -5
rect 389 -6 390 -5
rect 390 -6 391 -5
rect 391 -6 392 -5
rect 392 -6 393 -5
rect 393 -6 394 -5
rect 394 -6 395 -5
rect 395 -6 396 -5
rect 396 -6 397 -5
rect 397 -6 398 -5
rect 398 -6 399 -5
rect 399 -6 400 -5
rect 400 -6 401 -5
rect 401 -6 402 -5
rect 402 -6 403 -5
rect 403 -6 404 -5
rect 404 -6 405 -5
rect 405 -6 406 -5
rect 406 -6 407 -5
rect 407 -6 408 -5
rect 408 -6 409 -5
rect 409 -6 410 -5
rect 410 -6 411 -5
rect 411 -6 412 -5
rect 412 -6 413 -5
rect 413 -6 414 -5
rect 414 -6 415 -5
rect 415 -6 416 -5
rect 416 -6 417 -5
rect 417 -6 418 -5
rect 418 -6 419 -5
rect 419 -6 420 -5
rect 420 -6 421 -5
rect 421 -6 422 -5
rect 422 -6 423 -5
rect 423 -6 424 -5
rect 424 -6 425 -5
rect 425 -6 426 -5
rect 426 -6 427 -5
rect 427 -6 428 -5
rect 428 -6 429 -5
rect 429 -6 430 -5
rect 430 -6 431 -5
rect 431 -6 432 -5
rect 432 -6 433 -5
rect 433 -6 434 -5
rect 434 -6 435 -5
rect 435 -6 436 -5
rect 436 -6 437 -5
rect 437 -6 438 -5
rect 438 -6 439 -5
rect 439 -6 440 -5
rect 440 -6 441 -5
rect 441 -6 442 -5
rect 442 -6 443 -5
rect 443 -6 444 -5
rect 444 -6 445 -5
rect 445 -6 446 -5
rect 446 -6 447 -5
rect 447 -6 448 -5
rect 448 -6 449 -5
rect 449 -6 450 -5
rect 450 -6 451 -5
rect 451 -6 452 -5
rect 452 -6 453 -5
rect 453 -6 454 -5
rect 454 -6 455 -5
rect 455 -6 456 -5
rect 456 -6 457 -5
rect 457 -6 458 -5
rect 458 -6 459 -5
rect 459 -6 460 -5
rect 460 -6 461 -5
rect 461 -6 462 -5
rect 462 -6 463 -5
rect 463 -6 464 -5
rect 464 -6 465 -5
rect 465 -6 466 -5
rect 466 -6 467 -5
rect 467 -6 468 -5
rect 468 -6 469 -5
rect 469 -6 470 -5
rect 470 -6 471 -5
rect 471 -6 472 -5
rect 472 -6 473 -5
rect 473 -6 474 -5
rect 474 -6 475 -5
rect 475 -6 476 -5
rect 476 -6 477 -5
rect 477 -6 478 -5
rect 478 -6 479 -5
rect 479 -6 480 -5
rect 2 -7 3 -6
rect 3 -7 4 -6
rect 4 -7 5 -6
rect 5 -7 6 -6
rect 6 -7 7 -6
rect 7 -7 8 -6
rect 8 -7 9 -6
rect 9 -7 10 -6
rect 10 -7 11 -6
rect 11 -7 12 -6
rect 12 -7 13 -6
rect 13 -7 14 -6
rect 14 -7 15 -6
rect 18 -7 19 -6
rect 19 -7 20 -6
rect 20 -7 21 -6
rect 21 -7 22 -6
rect 22 -7 23 -6
rect 23 -7 24 -6
rect 24 -7 25 -6
rect 25 -7 26 -6
rect 26 -7 27 -6
rect 27 -7 28 -6
rect 28 -7 29 -6
rect 29 -7 30 -6
rect 30 -7 31 -6
rect 31 -7 32 -6
rect 32 -7 33 -6
rect 33 -7 34 -6
rect 34 -7 35 -6
rect 35 -7 36 -6
rect 36 -7 37 -6
rect 37 -7 38 -6
rect 38 -7 39 -6
rect 39 -7 40 -6
rect 40 -7 41 -6
rect 41 -7 42 -6
rect 42 -7 43 -6
rect 43 -7 44 -6
rect 44 -7 45 -6
rect 45 -7 46 -6
rect 46 -7 47 -6
rect 50 -7 51 -6
rect 51 -7 52 -6
rect 52 -7 53 -6
rect 53 -7 54 -6
rect 54 -7 55 -6
rect 55 -7 56 -6
rect 56 -7 57 -6
rect 57 -7 58 -6
rect 58 -7 59 -6
rect 59 -7 60 -6
rect 60 -7 61 -6
rect 61 -7 62 -6
rect 62 -7 63 -6
rect 63 -7 64 -6
rect 64 -7 65 -6
rect 65 -7 66 -6
rect 66 -7 67 -6
rect 67 -7 68 -6
rect 68 -7 69 -6
rect 69 -7 70 -6
rect 70 -7 71 -6
rect 71 -7 72 -6
rect 72 -7 73 -6
rect 73 -7 74 -6
rect 74 -7 75 -6
rect 75 -7 76 -6
rect 76 -7 77 -6
rect 77 -7 78 -6
rect 78 -7 79 -6
rect 82 -7 83 -6
rect 83 -7 84 -6
rect 84 -7 85 -6
rect 85 -7 86 -6
rect 86 -7 87 -6
rect 87 -7 88 -6
rect 88 -7 89 -6
rect 89 -7 90 -6
rect 90 -7 91 -6
rect 91 -7 92 -6
rect 92 -7 93 -6
rect 93 -7 94 -6
rect 94 -7 95 -6
rect 95 -7 96 -6
rect 96 -7 97 -6
rect 97 -7 98 -6
rect 98 -7 99 -6
rect 99 -7 100 -6
rect 100 -7 101 -6
rect 101 -7 102 -6
rect 102 -7 103 -6
rect 103 -7 104 -6
rect 104 -7 105 -6
rect 105 -7 106 -6
rect 106 -7 107 -6
rect 107 -7 108 -6
rect 108 -7 109 -6
rect 109 -7 110 -6
rect 110 -7 111 -6
rect 114 -7 115 -6
rect 115 -7 116 -6
rect 116 -7 117 -6
rect 117 -7 118 -6
rect 118 -7 119 -6
rect 119 -7 120 -6
rect 120 -7 121 -6
rect 121 -7 122 -6
rect 122 -7 123 -6
rect 123 -7 124 -6
rect 124 -7 125 -6
rect 125 -7 126 -6
rect 126 -7 127 -6
rect 127 -7 128 -6
rect 128 -7 129 -6
rect 129 -7 130 -6
rect 130 -7 131 -6
rect 131 -7 132 -6
rect 132 -7 133 -6
rect 133 -7 134 -6
rect 134 -7 135 -6
rect 135 -7 136 -6
rect 136 -7 137 -6
rect 137 -7 138 -6
rect 138 -7 139 -6
rect 139 -7 140 -6
rect 140 -7 141 -6
rect 141 -7 142 -6
rect 142 -7 143 -6
rect 146 -7 147 -6
rect 147 -7 148 -6
rect 148 -7 149 -6
rect 149 -7 150 -6
rect 150 -7 151 -6
rect 151 -7 152 -6
rect 152 -7 153 -6
rect 153 -7 154 -6
rect 154 -7 155 -6
rect 155 -7 156 -6
rect 156 -7 157 -6
rect 157 -7 158 -6
rect 158 -7 159 -6
rect 159 -7 160 -6
rect 160 -7 161 -6
rect 161 -7 162 -6
rect 162 -7 163 -6
rect 163 -7 164 -6
rect 164 -7 165 -6
rect 165 -7 166 -6
rect 166 -7 167 -6
rect 167 -7 168 -6
rect 168 -7 169 -6
rect 169 -7 170 -6
rect 170 -7 171 -6
rect 171 -7 172 -6
rect 172 -7 173 -6
rect 173 -7 174 -6
rect 174 -7 175 -6
rect 178 -7 179 -6
rect 179 -7 180 -6
rect 180 -7 181 -6
rect 181 -7 182 -6
rect 182 -7 183 -6
rect 183 -7 184 -6
rect 184 -7 185 -6
rect 185 -7 186 -6
rect 186 -7 187 -6
rect 187 -7 188 -6
rect 188 -7 189 -6
rect 189 -7 190 -6
rect 190 -7 191 -6
rect 191 -7 192 -6
rect 192 -7 193 -6
rect 193 -7 194 -6
rect 194 -7 195 -6
rect 195 -7 196 -6
rect 196 -7 197 -6
rect 197 -7 198 -6
rect 198 -7 199 -6
rect 199 -7 200 -6
rect 200 -7 201 -6
rect 201 -7 202 -6
rect 202 -7 203 -6
rect 203 -7 204 -6
rect 204 -7 205 -6
rect 205 -7 206 -6
rect 206 -7 207 -6
rect 207 -7 208 -6
rect 208 -7 209 -6
rect 209 -7 210 -6
rect 210 -7 211 -6
rect 211 -7 212 -6
rect 212 -7 213 -6
rect 213 -7 214 -6
rect 214 -7 215 -6
rect 215 -7 216 -6
rect 216 -7 217 -6
rect 217 -7 218 -6
rect 218 -7 219 -6
rect 219 -7 220 -6
rect 220 -7 221 -6
rect 221 -7 222 -6
rect 222 -7 223 -6
rect 223 -7 224 -6
rect 224 -7 225 -6
rect 225 -7 226 -6
rect 226 -7 227 -6
rect 227 -7 228 -6
rect 228 -7 229 -6
rect 229 -7 230 -6
rect 230 -7 231 -6
rect 231 -7 232 -6
rect 232 -7 233 -6
rect 233 -7 234 -6
rect 234 -7 235 -6
rect 235 -7 236 -6
rect 236 -7 237 -6
rect 237 -7 238 -6
rect 238 -7 239 -6
rect 239 -7 240 -6
rect 240 -7 241 -6
rect 241 -7 242 -6
rect 242 -7 243 -6
rect 243 -7 244 -6
rect 244 -7 245 -6
rect 245 -7 246 -6
rect 246 -7 247 -6
rect 247 -7 248 -6
rect 248 -7 249 -6
rect 249 -7 250 -6
rect 250 -7 251 -6
rect 251 -7 252 -6
rect 252 -7 253 -6
rect 253 -7 254 -6
rect 254 -7 255 -6
rect 255 -7 256 -6
rect 256 -7 257 -6
rect 257 -7 258 -6
rect 258 -7 259 -6
rect 259 -7 260 -6
rect 260 -7 261 -6
rect 261 -7 262 -6
rect 262 -7 263 -6
rect 263 -7 264 -6
rect 264 -7 265 -6
rect 265 -7 266 -6
rect 266 -7 267 -6
rect 267 -7 268 -6
rect 268 -7 269 -6
rect 269 -7 270 -6
rect 270 -7 271 -6
rect 271 -7 272 -6
rect 272 -7 273 -6
rect 273 -7 274 -6
rect 274 -7 275 -6
rect 275 -7 276 -6
rect 276 -7 277 -6
rect 277 -7 278 -6
rect 278 -7 279 -6
rect 279 -7 280 -6
rect 280 -7 281 -6
rect 281 -7 282 -6
rect 282 -7 283 -6
rect 283 -7 284 -6
rect 284 -7 285 -6
rect 285 -7 286 -6
rect 286 -7 287 -6
rect 287 -7 288 -6
rect 288 -7 289 -6
rect 289 -7 290 -6
rect 290 -7 291 -6
rect 291 -7 292 -6
rect 292 -7 293 -6
rect 293 -7 294 -6
rect 294 -7 295 -6
rect 295 -7 296 -6
rect 296 -7 297 -6
rect 297 -7 298 -6
rect 298 -7 299 -6
rect 299 -7 300 -6
rect 300 -7 301 -6
rect 301 -7 302 -6
rect 302 -7 303 -6
rect 303 -7 304 -6
rect 304 -7 305 -6
rect 305 -7 306 -6
rect 306 -7 307 -6
rect 307 -7 308 -6
rect 308 -7 309 -6
rect 309 -7 310 -6
rect 310 -7 311 -6
rect 311 -7 312 -6
rect 312 -7 313 -6
rect 313 -7 314 -6
rect 314 -7 315 -6
rect 315 -7 316 -6
rect 316 -7 317 -6
rect 317 -7 318 -6
rect 318 -7 319 -6
rect 319 -7 320 -6
rect 320 -7 321 -6
rect 321 -7 322 -6
rect 322 -7 323 -6
rect 323 -7 324 -6
rect 324 -7 325 -6
rect 325 -7 326 -6
rect 326 -7 327 -6
rect 327 -7 328 -6
rect 328 -7 329 -6
rect 329 -7 330 -6
rect 330 -7 331 -6
rect 331 -7 332 -6
rect 332 -7 333 -6
rect 333 -7 334 -6
rect 334 -7 335 -6
rect 335 -7 336 -6
rect 336 -7 337 -6
rect 337 -7 338 -6
rect 338 -7 339 -6
rect 339 -7 340 -6
rect 340 -7 341 -6
rect 341 -7 342 -6
rect 342 -7 343 -6
rect 343 -7 344 -6
rect 344 -7 345 -6
rect 345 -7 346 -6
rect 346 -7 347 -6
rect 347 -7 348 -6
rect 348 -7 349 -6
rect 349 -7 350 -6
rect 350 -7 351 -6
rect 351 -7 352 -6
rect 352 -7 353 -6
rect 353 -7 354 -6
rect 354 -7 355 -6
rect 355 -7 356 -6
rect 356 -7 357 -6
rect 357 -7 358 -6
rect 358 -7 359 -6
rect 359 -7 360 -6
rect 360 -7 361 -6
rect 361 -7 362 -6
rect 362 -7 363 -6
rect 363 -7 364 -6
rect 364 -7 365 -6
rect 365 -7 366 -6
rect 366 -7 367 -6
rect 367 -7 368 -6
rect 368 -7 369 -6
rect 369 -7 370 -6
rect 370 -7 371 -6
rect 371 -7 372 -6
rect 372 -7 373 -6
rect 373 -7 374 -6
rect 374 -7 375 -6
rect 375 -7 376 -6
rect 376 -7 377 -6
rect 377 -7 378 -6
rect 378 -7 379 -6
rect 379 -7 380 -6
rect 380 -7 381 -6
rect 381 -7 382 -6
rect 382 -7 383 -6
rect 383 -7 384 -6
rect 384 -7 385 -6
rect 385 -7 386 -6
rect 386 -7 387 -6
rect 387 -7 388 -6
rect 388 -7 389 -6
rect 389 -7 390 -6
rect 390 -7 391 -6
rect 391 -7 392 -6
rect 392 -7 393 -6
rect 393 -7 394 -6
rect 394 -7 395 -6
rect 395 -7 396 -6
rect 396 -7 397 -6
rect 397 -7 398 -6
rect 398 -7 399 -6
rect 399 -7 400 -6
rect 400 -7 401 -6
rect 401 -7 402 -6
rect 402 -7 403 -6
rect 403 -7 404 -6
rect 404 -7 405 -6
rect 405 -7 406 -6
rect 406 -7 407 -6
rect 407 -7 408 -6
rect 408 -7 409 -6
rect 409 -7 410 -6
rect 410 -7 411 -6
rect 411 -7 412 -6
rect 412 -7 413 -6
rect 413 -7 414 -6
rect 414 -7 415 -6
rect 415 -7 416 -6
rect 416 -7 417 -6
rect 417 -7 418 -6
rect 418 -7 419 -6
rect 419 -7 420 -6
rect 420 -7 421 -6
rect 421 -7 422 -6
rect 422 -7 423 -6
rect 423 -7 424 -6
rect 424 -7 425 -6
rect 425 -7 426 -6
rect 426 -7 427 -6
rect 427 -7 428 -6
rect 428 -7 429 -6
rect 429 -7 430 -6
rect 430 -7 431 -6
rect 431 -7 432 -6
rect 432 -7 433 -6
rect 433 -7 434 -6
rect 434 -7 435 -6
rect 435 -7 436 -6
rect 436 -7 437 -6
rect 437 -7 438 -6
rect 438 -7 439 -6
rect 439 -7 440 -6
rect 440 -7 441 -6
rect 441 -7 442 -6
rect 442 -7 443 -6
rect 443 -7 444 -6
rect 444 -7 445 -6
rect 445 -7 446 -6
rect 446 -7 447 -6
rect 447 -7 448 -6
rect 448 -7 449 -6
rect 449 -7 450 -6
rect 450 -7 451 -6
rect 451 -7 452 -6
rect 452 -7 453 -6
rect 453 -7 454 -6
rect 454 -7 455 -6
rect 455 -7 456 -6
rect 456 -7 457 -6
rect 457 -7 458 -6
rect 458 -7 459 -6
rect 459 -7 460 -6
rect 460 -7 461 -6
rect 461 -7 462 -6
rect 462 -7 463 -6
rect 463 -7 464 -6
rect 464 -7 465 -6
rect 465 -7 466 -6
rect 466 -7 467 -6
rect 467 -7 468 -6
rect 468 -7 469 -6
rect 469 -7 470 -6
rect 470 -7 471 -6
rect 471 -7 472 -6
rect 472 -7 473 -6
rect 473 -7 474 -6
rect 474 -7 475 -6
rect 475 -7 476 -6
rect 476 -7 477 -6
rect 477 -7 478 -6
rect 478 -7 479 -6
rect 479 -7 480 -6
rect 2 -8 3 -7
rect 3 -8 4 -7
rect 4 -8 5 -7
rect 5 -8 6 -7
rect 6 -8 7 -7
rect 7 -8 8 -7
rect 8 -8 9 -7
rect 9 -8 10 -7
rect 10 -8 11 -7
rect 11 -8 12 -7
rect 12 -8 13 -7
rect 13 -8 14 -7
rect 14 -8 15 -7
rect 19 -8 20 -7
rect 20 -8 21 -7
rect 21 -8 22 -7
rect 22 -8 23 -7
rect 23 -8 24 -7
rect 24 -8 25 -7
rect 25 -8 26 -7
rect 26 -8 27 -7
rect 27 -8 28 -7
rect 28 -8 29 -7
rect 29 -8 30 -7
rect 30 -8 31 -7
rect 31 -8 32 -7
rect 32 -8 33 -7
rect 33 -8 34 -7
rect 34 -8 35 -7
rect 35 -8 36 -7
rect 36 -8 37 -7
rect 37 -8 38 -7
rect 38 -8 39 -7
rect 39 -8 40 -7
rect 40 -8 41 -7
rect 41 -8 42 -7
rect 42 -8 43 -7
rect 43 -8 44 -7
rect 44 -8 45 -7
rect 45 -8 46 -7
rect 46 -8 47 -7
rect 51 -8 52 -7
rect 52 -8 53 -7
rect 53 -8 54 -7
rect 54 -8 55 -7
rect 55 -8 56 -7
rect 56 -8 57 -7
rect 57 -8 58 -7
rect 58 -8 59 -7
rect 59 -8 60 -7
rect 60 -8 61 -7
rect 61 -8 62 -7
rect 62 -8 63 -7
rect 63 -8 64 -7
rect 64 -8 65 -7
rect 65 -8 66 -7
rect 66 -8 67 -7
rect 67 -8 68 -7
rect 68 -8 69 -7
rect 69 -8 70 -7
rect 70 -8 71 -7
rect 71 -8 72 -7
rect 72 -8 73 -7
rect 73 -8 74 -7
rect 74 -8 75 -7
rect 75 -8 76 -7
rect 76 -8 77 -7
rect 77 -8 78 -7
rect 78 -8 79 -7
rect 83 -8 84 -7
rect 84 -8 85 -7
rect 85 -8 86 -7
rect 86 -8 87 -7
rect 87 -8 88 -7
rect 88 -8 89 -7
rect 89 -8 90 -7
rect 90 -8 91 -7
rect 91 -8 92 -7
rect 92 -8 93 -7
rect 93 -8 94 -7
rect 94 -8 95 -7
rect 95 -8 96 -7
rect 96 -8 97 -7
rect 97 -8 98 -7
rect 98 -8 99 -7
rect 99 -8 100 -7
rect 100 -8 101 -7
rect 101 -8 102 -7
rect 102 -8 103 -7
rect 103 -8 104 -7
rect 104 -8 105 -7
rect 105 -8 106 -7
rect 106 -8 107 -7
rect 107 -8 108 -7
rect 108 -8 109 -7
rect 109 -8 110 -7
rect 110 -8 111 -7
rect 115 -8 116 -7
rect 116 -8 117 -7
rect 117 -8 118 -7
rect 118 -8 119 -7
rect 119 -8 120 -7
rect 120 -8 121 -7
rect 121 -8 122 -7
rect 122 -8 123 -7
rect 123 -8 124 -7
rect 124 -8 125 -7
rect 125 -8 126 -7
rect 126 -8 127 -7
rect 127 -8 128 -7
rect 128 -8 129 -7
rect 129 -8 130 -7
rect 130 -8 131 -7
rect 131 -8 132 -7
rect 132 -8 133 -7
rect 133 -8 134 -7
rect 134 -8 135 -7
rect 135 -8 136 -7
rect 136 -8 137 -7
rect 137 -8 138 -7
rect 138 -8 139 -7
rect 139 -8 140 -7
rect 140 -8 141 -7
rect 141 -8 142 -7
rect 142 -8 143 -7
rect 147 -8 148 -7
rect 148 -8 149 -7
rect 149 -8 150 -7
rect 150 -8 151 -7
rect 151 -8 152 -7
rect 152 -8 153 -7
rect 153 -8 154 -7
rect 154 -8 155 -7
rect 155 -8 156 -7
rect 156 -8 157 -7
rect 157 -8 158 -7
rect 158 -8 159 -7
rect 159 -8 160 -7
rect 160 -8 161 -7
rect 161 -8 162 -7
rect 162 -8 163 -7
rect 163 -8 164 -7
rect 164 -8 165 -7
rect 165 -8 166 -7
rect 166 -8 167 -7
rect 167 -8 168 -7
rect 168 -8 169 -7
rect 169 -8 170 -7
rect 170 -8 171 -7
rect 171 -8 172 -7
rect 172 -8 173 -7
rect 173 -8 174 -7
rect 174 -8 175 -7
rect 179 -8 180 -7
rect 180 -8 181 -7
rect 181 -8 182 -7
rect 182 -8 183 -7
rect 183 -8 184 -7
rect 184 -8 185 -7
rect 185 -8 186 -7
rect 186 -8 187 -7
rect 187 -8 188 -7
rect 188 -8 189 -7
rect 189 -8 190 -7
rect 190 -8 191 -7
rect 191 -8 192 -7
rect 192 -8 193 -7
rect 193 -8 194 -7
rect 194 -8 195 -7
rect 195 -8 196 -7
rect 196 -8 197 -7
rect 197 -8 198 -7
rect 198 -8 199 -7
rect 199 -8 200 -7
rect 200 -8 201 -7
rect 201 -8 202 -7
rect 202 -8 203 -7
rect 203 -8 204 -7
rect 204 -8 205 -7
rect 205 -8 206 -7
rect 206 -8 207 -7
rect 207 -8 208 -7
rect 208 -8 209 -7
rect 209 -8 210 -7
rect 210 -8 211 -7
rect 211 -8 212 -7
rect 212 -8 213 -7
rect 213 -8 214 -7
rect 214 -8 215 -7
rect 215 -8 216 -7
rect 216 -8 217 -7
rect 217 -8 218 -7
rect 218 -8 219 -7
rect 219 -8 220 -7
rect 220 -8 221 -7
rect 221 -8 222 -7
rect 222 -8 223 -7
rect 223 -8 224 -7
rect 224 -8 225 -7
rect 225 -8 226 -7
rect 226 -8 227 -7
rect 227 -8 228 -7
rect 228 -8 229 -7
rect 229 -8 230 -7
rect 230 -8 231 -7
rect 231 -8 232 -7
rect 232 -8 233 -7
rect 233 -8 234 -7
rect 234 -8 235 -7
rect 235 -8 236 -7
rect 236 -8 237 -7
rect 237 -8 238 -7
rect 238 -8 239 -7
rect 239 -8 240 -7
rect 240 -8 241 -7
rect 241 -8 242 -7
rect 242 -8 243 -7
rect 243 -8 244 -7
rect 244 -8 245 -7
rect 245 -8 246 -7
rect 246 -8 247 -7
rect 247 -8 248 -7
rect 248 -8 249 -7
rect 249 -8 250 -7
rect 250 -8 251 -7
rect 251 -8 252 -7
rect 252 -8 253 -7
rect 253 -8 254 -7
rect 254 -8 255 -7
rect 255 -8 256 -7
rect 256 -8 257 -7
rect 257 -8 258 -7
rect 258 -8 259 -7
rect 259 -8 260 -7
rect 260 -8 261 -7
rect 261 -8 262 -7
rect 262 -8 263 -7
rect 263 -8 264 -7
rect 264 -8 265 -7
rect 265 -8 266 -7
rect 266 -8 267 -7
rect 267 -8 268 -7
rect 268 -8 269 -7
rect 269 -8 270 -7
rect 270 -8 271 -7
rect 271 -8 272 -7
rect 272 -8 273 -7
rect 273 -8 274 -7
rect 274 -8 275 -7
rect 275 -8 276 -7
rect 276 -8 277 -7
rect 277 -8 278 -7
rect 278 -8 279 -7
rect 279 -8 280 -7
rect 280 -8 281 -7
rect 281 -8 282 -7
rect 282 -8 283 -7
rect 283 -8 284 -7
rect 284 -8 285 -7
rect 285 -8 286 -7
rect 286 -8 287 -7
rect 287 -8 288 -7
rect 288 -8 289 -7
rect 289 -8 290 -7
rect 290 -8 291 -7
rect 291 -8 292 -7
rect 292 -8 293 -7
rect 293 -8 294 -7
rect 294 -8 295 -7
rect 295 -8 296 -7
rect 296 -8 297 -7
rect 297 -8 298 -7
rect 298 -8 299 -7
rect 299 -8 300 -7
rect 300 -8 301 -7
rect 301 -8 302 -7
rect 302 -8 303 -7
rect 303 -8 304 -7
rect 304 -8 305 -7
rect 305 -8 306 -7
rect 306 -8 307 -7
rect 307 -8 308 -7
rect 308 -8 309 -7
rect 309 -8 310 -7
rect 310 -8 311 -7
rect 311 -8 312 -7
rect 312 -8 313 -7
rect 313 -8 314 -7
rect 314 -8 315 -7
rect 315 -8 316 -7
rect 316 -8 317 -7
rect 317 -8 318 -7
rect 318 -8 319 -7
rect 319 -8 320 -7
rect 320 -8 321 -7
rect 321 -8 322 -7
rect 322 -8 323 -7
rect 323 -8 324 -7
rect 324 -8 325 -7
rect 325 -8 326 -7
rect 326 -8 327 -7
rect 327 -8 328 -7
rect 328 -8 329 -7
rect 329 -8 330 -7
rect 330 -8 331 -7
rect 331 -8 332 -7
rect 332 -8 333 -7
rect 333 -8 334 -7
rect 334 -8 335 -7
rect 335 -8 336 -7
rect 336 -8 337 -7
rect 337 -8 338 -7
rect 338 -8 339 -7
rect 339 -8 340 -7
rect 340 -8 341 -7
rect 341 -8 342 -7
rect 342 -8 343 -7
rect 343 -8 344 -7
rect 344 -8 345 -7
rect 345 -8 346 -7
rect 346 -8 347 -7
rect 347 -8 348 -7
rect 348 -8 349 -7
rect 349 -8 350 -7
rect 350 -8 351 -7
rect 351 -8 352 -7
rect 352 -8 353 -7
rect 353 -8 354 -7
rect 354 -8 355 -7
rect 355 -8 356 -7
rect 356 -8 357 -7
rect 357 -8 358 -7
rect 358 -8 359 -7
rect 359 -8 360 -7
rect 360 -8 361 -7
rect 361 -8 362 -7
rect 362 -8 363 -7
rect 363 -8 364 -7
rect 364 -8 365 -7
rect 365 -8 366 -7
rect 366 -8 367 -7
rect 367 -8 368 -7
rect 368 -8 369 -7
rect 369 -8 370 -7
rect 370 -8 371 -7
rect 371 -8 372 -7
rect 372 -8 373 -7
rect 373 -8 374 -7
rect 374 -8 375 -7
rect 375 -8 376 -7
rect 376 -8 377 -7
rect 377 -8 378 -7
rect 378 -8 379 -7
rect 379 -8 380 -7
rect 380 -8 381 -7
rect 381 -8 382 -7
rect 382 -8 383 -7
rect 383 -8 384 -7
rect 384 -8 385 -7
rect 385 -8 386 -7
rect 386 -8 387 -7
rect 387 -8 388 -7
rect 388 -8 389 -7
rect 389 -8 390 -7
rect 390 -8 391 -7
rect 391 -8 392 -7
rect 392 -8 393 -7
rect 393 -8 394 -7
rect 394 -8 395 -7
rect 395 -8 396 -7
rect 396 -8 397 -7
rect 397 -8 398 -7
rect 398 -8 399 -7
rect 399 -8 400 -7
rect 400 -8 401 -7
rect 401 -8 402 -7
rect 402 -8 403 -7
rect 403 -8 404 -7
rect 404 -8 405 -7
rect 405 -8 406 -7
rect 406 -8 407 -7
rect 407 -8 408 -7
rect 408 -8 409 -7
rect 409 -8 410 -7
rect 410 -8 411 -7
rect 411 -8 412 -7
rect 412 -8 413 -7
rect 413 -8 414 -7
rect 414 -8 415 -7
rect 415 -8 416 -7
rect 416 -8 417 -7
rect 417 -8 418 -7
rect 418 -8 419 -7
rect 419 -8 420 -7
rect 420 -8 421 -7
rect 421 -8 422 -7
rect 422 -8 423 -7
rect 423 -8 424 -7
rect 424 -8 425 -7
rect 425 -8 426 -7
rect 426 -8 427 -7
rect 427 -8 428 -7
rect 428 -8 429 -7
rect 429 -8 430 -7
rect 430 -8 431 -7
rect 431 -8 432 -7
rect 432 -8 433 -7
rect 433 -8 434 -7
rect 434 -8 435 -7
rect 435 -8 436 -7
rect 436 -8 437 -7
rect 437 -8 438 -7
rect 438 -8 439 -7
rect 439 -8 440 -7
rect 440 -8 441 -7
rect 441 -8 442 -7
rect 442 -8 443 -7
rect 443 -8 444 -7
rect 444 -8 445 -7
rect 445 -8 446 -7
rect 446 -8 447 -7
rect 447 -8 448 -7
rect 448 -8 449 -7
rect 449 -8 450 -7
rect 450 -8 451 -7
rect 451 -8 452 -7
rect 452 -8 453 -7
rect 453 -8 454 -7
rect 454 -8 455 -7
rect 455 -8 456 -7
rect 456 -8 457 -7
rect 457 -8 458 -7
rect 458 -8 459 -7
rect 459 -8 460 -7
rect 460 -8 461 -7
rect 461 -8 462 -7
rect 462 -8 463 -7
rect 463 -8 464 -7
rect 464 -8 465 -7
rect 465 -8 466 -7
rect 466 -8 467 -7
rect 467 -8 468 -7
rect 468 -8 469 -7
rect 469 -8 470 -7
rect 470 -8 471 -7
rect 471 -8 472 -7
rect 472 -8 473 -7
rect 473 -8 474 -7
rect 474 -8 475 -7
rect 475 -8 476 -7
rect 476 -8 477 -7
rect 477 -8 478 -7
rect 478 -8 479 -7
rect 479 -8 480 -7
rect 2 -9 3 -8
rect 3 -9 4 -8
rect 4 -9 5 -8
rect 5 -9 6 -8
rect 6 -9 7 -8
rect 7 -9 8 -8
rect 8 -9 9 -8
rect 9 -9 10 -8
rect 10 -9 11 -8
rect 11 -9 12 -8
rect 12 -9 13 -8
rect 13 -9 14 -8
rect 19 -9 20 -8
rect 20 -9 21 -8
rect 21 -9 22 -8
rect 22 -9 23 -8
rect 23 -9 24 -8
rect 24 -9 25 -8
rect 25 -9 26 -8
rect 26 -9 27 -8
rect 27 -9 28 -8
rect 28 -9 29 -8
rect 29 -9 30 -8
rect 30 -9 31 -8
rect 31 -9 32 -8
rect 32 -9 33 -8
rect 33 -9 34 -8
rect 34 -9 35 -8
rect 35 -9 36 -8
rect 36 -9 37 -8
rect 37 -9 38 -8
rect 38 -9 39 -8
rect 39 -9 40 -8
rect 40 -9 41 -8
rect 41 -9 42 -8
rect 42 -9 43 -8
rect 43 -9 44 -8
rect 44 -9 45 -8
rect 45 -9 46 -8
rect 51 -9 52 -8
rect 52 -9 53 -8
rect 53 -9 54 -8
rect 54 -9 55 -8
rect 55 -9 56 -8
rect 56 -9 57 -8
rect 57 -9 58 -8
rect 58 -9 59 -8
rect 59 -9 60 -8
rect 60 -9 61 -8
rect 61 -9 62 -8
rect 62 -9 63 -8
rect 63 -9 64 -8
rect 64 -9 65 -8
rect 65 -9 66 -8
rect 66 -9 67 -8
rect 67 -9 68 -8
rect 68 -9 69 -8
rect 69 -9 70 -8
rect 70 -9 71 -8
rect 71 -9 72 -8
rect 72 -9 73 -8
rect 73 -9 74 -8
rect 74 -9 75 -8
rect 75 -9 76 -8
rect 76 -9 77 -8
rect 77 -9 78 -8
rect 83 -9 84 -8
rect 84 -9 85 -8
rect 85 -9 86 -8
rect 86 -9 87 -8
rect 87 -9 88 -8
rect 88 -9 89 -8
rect 89 -9 90 -8
rect 90 -9 91 -8
rect 91 -9 92 -8
rect 92 -9 93 -8
rect 93 -9 94 -8
rect 94 -9 95 -8
rect 95 -9 96 -8
rect 96 -9 97 -8
rect 97 -9 98 -8
rect 98 -9 99 -8
rect 99 -9 100 -8
rect 100 -9 101 -8
rect 101 -9 102 -8
rect 102 -9 103 -8
rect 103 -9 104 -8
rect 104 -9 105 -8
rect 105 -9 106 -8
rect 106 -9 107 -8
rect 107 -9 108 -8
rect 108 -9 109 -8
rect 109 -9 110 -8
rect 115 -9 116 -8
rect 116 -9 117 -8
rect 117 -9 118 -8
rect 118 -9 119 -8
rect 119 -9 120 -8
rect 120 -9 121 -8
rect 121 -9 122 -8
rect 122 -9 123 -8
rect 123 -9 124 -8
rect 124 -9 125 -8
rect 125 -9 126 -8
rect 126 -9 127 -8
rect 127 -9 128 -8
rect 128 -9 129 -8
rect 129 -9 130 -8
rect 130 -9 131 -8
rect 131 -9 132 -8
rect 132 -9 133 -8
rect 133 -9 134 -8
rect 134 -9 135 -8
rect 135 -9 136 -8
rect 136 -9 137 -8
rect 137 -9 138 -8
rect 138 -9 139 -8
rect 139 -9 140 -8
rect 140 -9 141 -8
rect 141 -9 142 -8
rect 147 -9 148 -8
rect 148 -9 149 -8
rect 149 -9 150 -8
rect 150 -9 151 -8
rect 151 -9 152 -8
rect 152 -9 153 -8
rect 153 -9 154 -8
rect 154 -9 155 -8
rect 155 -9 156 -8
rect 156 -9 157 -8
rect 157 -9 158 -8
rect 158 -9 159 -8
rect 159 -9 160 -8
rect 160 -9 161 -8
rect 161 -9 162 -8
rect 162 -9 163 -8
rect 163 -9 164 -8
rect 164 -9 165 -8
rect 165 -9 166 -8
rect 166 -9 167 -8
rect 167 -9 168 -8
rect 168 -9 169 -8
rect 169 -9 170 -8
rect 170 -9 171 -8
rect 171 -9 172 -8
rect 172 -9 173 -8
rect 173 -9 174 -8
rect 179 -9 180 -8
rect 180 -9 181 -8
rect 181 -9 182 -8
rect 182 -9 183 -8
rect 183 -9 184 -8
rect 184 -9 185 -8
rect 185 -9 186 -8
rect 186 -9 187 -8
rect 187 -9 188 -8
rect 188 -9 189 -8
rect 189 -9 190 -8
rect 190 -9 191 -8
rect 191 -9 192 -8
rect 192 -9 193 -8
rect 193 -9 194 -8
rect 194 -9 195 -8
rect 195 -9 196 -8
rect 196 -9 197 -8
rect 197 -9 198 -8
rect 198 -9 199 -8
rect 199 -9 200 -8
rect 200 -9 201 -8
rect 201 -9 202 -8
rect 202 -9 203 -8
rect 203 -9 204 -8
rect 204 -9 205 -8
rect 205 -9 206 -8
rect 206 -9 207 -8
rect 207 -9 208 -8
rect 208 -9 209 -8
rect 209 -9 210 -8
rect 210 -9 211 -8
rect 211 -9 212 -8
rect 212 -9 213 -8
rect 213 -9 214 -8
rect 214 -9 215 -8
rect 215 -9 216 -8
rect 216 -9 217 -8
rect 217 -9 218 -8
rect 218 -9 219 -8
rect 219 -9 220 -8
rect 220 -9 221 -8
rect 221 -9 222 -8
rect 222 -9 223 -8
rect 223 -9 224 -8
rect 224 -9 225 -8
rect 225 -9 226 -8
rect 226 -9 227 -8
rect 227 -9 228 -8
rect 228 -9 229 -8
rect 229 -9 230 -8
rect 230 -9 231 -8
rect 231 -9 232 -8
rect 232 -9 233 -8
rect 233 -9 234 -8
rect 234 -9 235 -8
rect 235 -9 236 -8
rect 236 -9 237 -8
rect 237 -9 238 -8
rect 238 -9 239 -8
rect 239 -9 240 -8
rect 240 -9 241 -8
rect 241 -9 242 -8
rect 242 -9 243 -8
rect 243 -9 244 -8
rect 244 -9 245 -8
rect 245 -9 246 -8
rect 246 -9 247 -8
rect 247 -9 248 -8
rect 248 -9 249 -8
rect 249 -9 250 -8
rect 250 -9 251 -8
rect 251 -9 252 -8
rect 252 -9 253 -8
rect 253 -9 254 -8
rect 254 -9 255 -8
rect 255 -9 256 -8
rect 256 -9 257 -8
rect 257 -9 258 -8
rect 258 -9 259 -8
rect 259 -9 260 -8
rect 260 -9 261 -8
rect 261 -9 262 -8
rect 262 -9 263 -8
rect 263 -9 264 -8
rect 264 -9 265 -8
rect 265 -9 266 -8
rect 266 -9 267 -8
rect 267 -9 268 -8
rect 268 -9 269 -8
rect 269 -9 270 -8
rect 270 -9 271 -8
rect 271 -9 272 -8
rect 272 -9 273 -8
rect 273 -9 274 -8
rect 274 -9 275 -8
rect 275 -9 276 -8
rect 276 -9 277 -8
rect 277 -9 278 -8
rect 278 -9 279 -8
rect 279 -9 280 -8
rect 280 -9 281 -8
rect 281 -9 282 -8
rect 282 -9 283 -8
rect 283 -9 284 -8
rect 284 -9 285 -8
rect 285 -9 286 -8
rect 286 -9 287 -8
rect 287 -9 288 -8
rect 288 -9 289 -8
rect 289 -9 290 -8
rect 290 -9 291 -8
rect 291 -9 292 -8
rect 292 -9 293 -8
rect 293 -9 294 -8
rect 294 -9 295 -8
rect 295 -9 296 -8
rect 296 -9 297 -8
rect 297 -9 298 -8
rect 298 -9 299 -8
rect 299 -9 300 -8
rect 300 -9 301 -8
rect 301 -9 302 -8
rect 302 -9 303 -8
rect 303 -9 304 -8
rect 304 -9 305 -8
rect 305 -9 306 -8
rect 306 -9 307 -8
rect 307 -9 308 -8
rect 308 -9 309 -8
rect 309 -9 310 -8
rect 310 -9 311 -8
rect 311 -9 312 -8
rect 312 -9 313 -8
rect 313 -9 314 -8
rect 314 -9 315 -8
rect 315 -9 316 -8
rect 316 -9 317 -8
rect 317 -9 318 -8
rect 318 -9 319 -8
rect 319 -9 320 -8
rect 320 -9 321 -8
rect 321 -9 322 -8
rect 322 -9 323 -8
rect 323 -9 324 -8
rect 324 -9 325 -8
rect 325 -9 326 -8
rect 326 -9 327 -8
rect 327 -9 328 -8
rect 328 -9 329 -8
rect 329 -9 330 -8
rect 330 -9 331 -8
rect 331 -9 332 -8
rect 332 -9 333 -8
rect 333 -9 334 -8
rect 334 -9 335 -8
rect 335 -9 336 -8
rect 336 -9 337 -8
rect 337 -9 338 -8
rect 338 -9 339 -8
rect 339 -9 340 -8
rect 340 -9 341 -8
rect 341 -9 342 -8
rect 342 -9 343 -8
rect 343 -9 344 -8
rect 344 -9 345 -8
rect 345 -9 346 -8
rect 346 -9 347 -8
rect 347 -9 348 -8
rect 348 -9 349 -8
rect 349 -9 350 -8
rect 350 -9 351 -8
rect 351 -9 352 -8
rect 352 -9 353 -8
rect 353 -9 354 -8
rect 354 -9 355 -8
rect 355 -9 356 -8
rect 356 -9 357 -8
rect 357 -9 358 -8
rect 358 -9 359 -8
rect 359 -9 360 -8
rect 360 -9 361 -8
rect 361 -9 362 -8
rect 362 -9 363 -8
rect 363 -9 364 -8
rect 364 -9 365 -8
rect 365 -9 366 -8
rect 366 -9 367 -8
rect 367 -9 368 -8
rect 368 -9 369 -8
rect 369 -9 370 -8
rect 370 -9 371 -8
rect 371 -9 372 -8
rect 372 -9 373 -8
rect 373 -9 374 -8
rect 374 -9 375 -8
rect 375 -9 376 -8
rect 376 -9 377 -8
rect 377 -9 378 -8
rect 378 -9 379 -8
rect 379 -9 380 -8
rect 380 -9 381 -8
rect 381 -9 382 -8
rect 382 -9 383 -8
rect 383 -9 384 -8
rect 384 -9 385 -8
rect 385 -9 386 -8
rect 386 -9 387 -8
rect 387 -9 388 -8
rect 388 -9 389 -8
rect 389 -9 390 -8
rect 390 -9 391 -8
rect 391 -9 392 -8
rect 392 -9 393 -8
rect 393 -9 394 -8
rect 394 -9 395 -8
rect 395 -9 396 -8
rect 396 -9 397 -8
rect 397 -9 398 -8
rect 398 -9 399 -8
rect 399 -9 400 -8
rect 400 -9 401 -8
rect 401 -9 402 -8
rect 402 -9 403 -8
rect 403 -9 404 -8
rect 404 -9 405 -8
rect 405 -9 406 -8
rect 406 -9 407 -8
rect 407 -9 408 -8
rect 408 -9 409 -8
rect 409 -9 410 -8
rect 410 -9 411 -8
rect 411 -9 412 -8
rect 412 -9 413 -8
rect 413 -9 414 -8
rect 414 -9 415 -8
rect 415 -9 416 -8
rect 416 -9 417 -8
rect 417 -9 418 -8
rect 418 -9 419 -8
rect 419 -9 420 -8
rect 420 -9 421 -8
rect 421 -9 422 -8
rect 422 -9 423 -8
rect 423 -9 424 -8
rect 424 -9 425 -8
rect 425 -9 426 -8
rect 426 -9 427 -8
rect 427 -9 428 -8
rect 428 -9 429 -8
rect 429 -9 430 -8
rect 430 -9 431 -8
rect 431 -9 432 -8
rect 432 -9 433 -8
rect 433 -9 434 -8
rect 434 -9 435 -8
rect 435 -9 436 -8
rect 436 -9 437 -8
rect 437 -9 438 -8
rect 438 -9 439 -8
rect 439 -9 440 -8
rect 440 -9 441 -8
rect 441 -9 442 -8
rect 442 -9 443 -8
rect 443 -9 444 -8
rect 444 -9 445 -8
rect 445 -9 446 -8
rect 446 -9 447 -8
rect 447 -9 448 -8
rect 448 -9 449 -8
rect 449 -9 450 -8
rect 450 -9 451 -8
rect 451 -9 452 -8
rect 452 -9 453 -8
rect 453 -9 454 -8
rect 454 -9 455 -8
rect 455 -9 456 -8
rect 456 -9 457 -8
rect 457 -9 458 -8
rect 458 -9 459 -8
rect 459 -9 460 -8
rect 460 -9 461 -8
rect 461 -9 462 -8
rect 462 -9 463 -8
rect 463 -9 464 -8
rect 464 -9 465 -8
rect 465 -9 466 -8
rect 466 -9 467 -8
rect 467 -9 468 -8
rect 468 -9 469 -8
rect 469 -9 470 -8
rect 470 -9 471 -8
rect 471 -9 472 -8
rect 472 -9 473 -8
rect 473 -9 474 -8
rect 474 -9 475 -8
rect 475 -9 476 -8
rect 476 -9 477 -8
rect 477 -9 478 -8
rect 478 -9 479 -8
rect 479 -9 480 -8
rect 2 -10 3 -9
rect 3 -10 4 -9
rect 4 -10 5 -9
rect 5 -10 6 -9
rect 6 -10 7 -9
rect 7 -10 8 -9
rect 8 -10 9 -9
rect 25 -10 26 -9
rect 26 -10 27 -9
rect 27 -10 28 -9
rect 28 -10 29 -9
rect 29 -10 30 -9
rect 30 -10 31 -9
rect 31 -10 32 -9
rect 32 -10 33 -9
rect 33 -10 34 -9
rect 34 -10 35 -9
rect 35 -10 36 -9
rect 36 -10 37 -9
rect 37 -10 38 -9
rect 38 -10 39 -9
rect 39 -10 40 -9
rect 40 -10 41 -9
rect 57 -10 58 -9
rect 58 -10 59 -9
rect 59 -10 60 -9
rect 60 -10 61 -9
rect 61 -10 62 -9
rect 62 -10 63 -9
rect 63 -10 64 -9
rect 64 -10 65 -9
rect 65 -10 66 -9
rect 66 -10 67 -9
rect 67 -10 68 -9
rect 68 -10 69 -9
rect 69 -10 70 -9
rect 70 -10 71 -9
rect 71 -10 72 -9
rect 72 -10 73 -9
rect 89 -10 90 -9
rect 90 -10 91 -9
rect 91 -10 92 -9
rect 92 -10 93 -9
rect 93 -10 94 -9
rect 94 -10 95 -9
rect 95 -10 96 -9
rect 96 -10 97 -9
rect 97 -10 98 -9
rect 98 -10 99 -9
rect 99 -10 100 -9
rect 100 -10 101 -9
rect 101 -10 102 -9
rect 102 -10 103 -9
rect 103 -10 104 -9
rect 104 -10 105 -9
rect 121 -10 122 -9
rect 122 -10 123 -9
rect 123 -10 124 -9
rect 124 -10 125 -9
rect 125 -10 126 -9
rect 126 -10 127 -9
rect 127 -10 128 -9
rect 128 -10 129 -9
rect 129 -10 130 -9
rect 130 -10 131 -9
rect 131 -10 132 -9
rect 132 -10 133 -9
rect 133 -10 134 -9
rect 134 -10 135 -9
rect 135 -10 136 -9
rect 136 -10 137 -9
rect 153 -10 154 -9
rect 154 -10 155 -9
rect 155 -10 156 -9
rect 156 -10 157 -9
rect 157 -10 158 -9
rect 158 -10 159 -9
rect 159 -10 160 -9
rect 160 -10 161 -9
rect 161 -10 162 -9
rect 162 -10 163 -9
rect 163 -10 164 -9
rect 164 -10 165 -9
rect 165 -10 166 -9
rect 166 -10 167 -9
rect 167 -10 168 -9
rect 168 -10 169 -9
rect 185 -10 186 -9
rect 186 -10 187 -9
rect 187 -10 188 -9
rect 188 -10 189 -9
rect 189 -10 190 -9
rect 190 -10 191 -9
rect 191 -10 192 -9
rect 192 -10 193 -9
rect 193 -10 194 -9
rect 194 -10 195 -9
rect 195 -10 196 -9
rect 196 -10 197 -9
rect 197 -10 198 -9
rect 198 -10 199 -9
rect 199 -10 200 -9
rect 200 -10 201 -9
rect 201 -10 202 -9
rect 202 -10 203 -9
rect 203 -10 204 -9
rect 204 -10 205 -9
rect 205 -10 206 -9
rect 206 -10 207 -9
rect 207 -10 208 -9
rect 208 -10 209 -9
rect 209 -10 210 -9
rect 210 -10 211 -9
rect 211 -10 212 -9
rect 212 -10 213 -9
rect 213 -10 214 -9
rect 214 -10 215 -9
rect 215 -10 216 -9
rect 216 -10 217 -9
rect 217 -10 218 -9
rect 218 -10 219 -9
rect 219 -10 220 -9
rect 220 -10 221 -9
rect 221 -10 222 -9
rect 222 -10 223 -9
rect 223 -10 224 -9
rect 224 -10 225 -9
rect 225 -10 226 -9
rect 226 -10 227 -9
rect 227 -10 228 -9
rect 228 -10 229 -9
rect 229 -10 230 -9
rect 230 -10 231 -9
rect 231 -10 232 -9
rect 232 -10 233 -9
rect 233 -10 234 -9
rect 234 -10 235 -9
rect 235 -10 236 -9
rect 236 -10 237 -9
rect 237 -10 238 -9
rect 238 -10 239 -9
rect 239 -10 240 -9
rect 240 -10 241 -9
rect 241 -10 242 -9
rect 242 -10 243 -9
rect 243 -10 244 -9
rect 244 -10 245 -9
rect 245 -10 246 -9
rect 246 -10 247 -9
rect 247 -10 248 -9
rect 248 -10 249 -9
rect 249 -10 250 -9
rect 250 -10 251 -9
rect 251 -10 252 -9
rect 252 -10 253 -9
rect 253 -10 254 -9
rect 254 -10 255 -9
rect 255 -10 256 -9
rect 256 -10 257 -9
rect 257 -10 258 -9
rect 258 -10 259 -9
rect 259 -10 260 -9
rect 260 -10 261 -9
rect 261 -10 262 -9
rect 262 -10 263 -9
rect 263 -10 264 -9
rect 264 -10 265 -9
rect 265 -10 266 -9
rect 266 -10 267 -9
rect 267 -10 268 -9
rect 268 -10 269 -9
rect 269 -10 270 -9
rect 270 -10 271 -9
rect 271 -10 272 -9
rect 272 -10 273 -9
rect 273 -10 274 -9
rect 274 -10 275 -9
rect 275 -10 276 -9
rect 276 -10 277 -9
rect 277 -10 278 -9
rect 278 -10 279 -9
rect 279 -10 280 -9
rect 280 -10 281 -9
rect 281 -10 282 -9
rect 282 -10 283 -9
rect 283 -10 284 -9
rect 284 -10 285 -9
rect 285 -10 286 -9
rect 286 -10 287 -9
rect 287 -10 288 -9
rect 288 -10 289 -9
rect 289 -10 290 -9
rect 290 -10 291 -9
rect 291 -10 292 -9
rect 292 -10 293 -9
rect 293 -10 294 -9
rect 294 -10 295 -9
rect 295 -10 296 -9
rect 296 -10 297 -9
rect 297 -10 298 -9
rect 298 -10 299 -9
rect 299 -10 300 -9
rect 300 -10 301 -9
rect 301 -10 302 -9
rect 302 -10 303 -9
rect 303 -10 304 -9
rect 304 -10 305 -9
rect 305 -10 306 -9
rect 306 -10 307 -9
rect 307 -10 308 -9
rect 308 -10 309 -9
rect 309 -10 310 -9
rect 310 -10 311 -9
rect 311 -10 312 -9
rect 312 -10 313 -9
rect 313 -10 314 -9
rect 314 -10 315 -9
rect 315 -10 316 -9
rect 316 -10 317 -9
rect 317 -10 318 -9
rect 318 -10 319 -9
rect 319 -10 320 -9
rect 320 -10 321 -9
rect 321 -10 322 -9
rect 322 -10 323 -9
rect 323 -10 324 -9
rect 324 -10 325 -9
rect 325 -10 326 -9
rect 326 -10 327 -9
rect 327 -10 328 -9
rect 328 -10 329 -9
rect 329 -10 330 -9
rect 330 -10 331 -9
rect 331 -10 332 -9
rect 332 -10 333 -9
rect 333 -10 334 -9
rect 334 -10 335 -9
rect 335 -10 336 -9
rect 336 -10 337 -9
rect 337 -10 338 -9
rect 338 -10 339 -9
rect 339 -10 340 -9
rect 340 -10 341 -9
rect 341 -10 342 -9
rect 342 -10 343 -9
rect 343 -10 344 -9
rect 344 -10 345 -9
rect 345 -10 346 -9
rect 346 -10 347 -9
rect 347 -10 348 -9
rect 348 -10 349 -9
rect 349 -10 350 -9
rect 350 -10 351 -9
rect 351 -10 352 -9
rect 352 -10 353 -9
rect 353 -10 354 -9
rect 354 -10 355 -9
rect 355 -10 356 -9
rect 356 -10 357 -9
rect 357 -10 358 -9
rect 358 -10 359 -9
rect 359 -10 360 -9
rect 360 -10 361 -9
rect 361 -10 362 -9
rect 362 -10 363 -9
rect 363 -10 364 -9
rect 364 -10 365 -9
rect 365 -10 366 -9
rect 366 -10 367 -9
rect 367 -10 368 -9
rect 368 -10 369 -9
rect 369 -10 370 -9
rect 370 -10 371 -9
rect 371 -10 372 -9
rect 372 -10 373 -9
rect 373 -10 374 -9
rect 374 -10 375 -9
rect 375 -10 376 -9
rect 376 -10 377 -9
rect 377 -10 378 -9
rect 378 -10 379 -9
rect 379 -10 380 -9
rect 380 -10 381 -9
rect 381 -10 382 -9
rect 382 -10 383 -9
rect 383 -10 384 -9
rect 384 -10 385 -9
rect 385 -10 386 -9
rect 386 -10 387 -9
rect 387 -10 388 -9
rect 388 -10 389 -9
rect 389 -10 390 -9
rect 390 -10 391 -9
rect 391 -10 392 -9
rect 392 -10 393 -9
rect 393 -10 394 -9
rect 394 -10 395 -9
rect 395 -10 396 -9
rect 396 -10 397 -9
rect 397 -10 398 -9
rect 398 -10 399 -9
rect 399 -10 400 -9
rect 400 -10 401 -9
rect 401 -10 402 -9
rect 402 -10 403 -9
rect 403 -10 404 -9
rect 404 -10 405 -9
rect 405 -10 406 -9
rect 406 -10 407 -9
rect 407 -10 408 -9
rect 408 -10 409 -9
rect 409 -10 410 -9
rect 410 -10 411 -9
rect 411 -10 412 -9
rect 412 -10 413 -9
rect 413 -10 414 -9
rect 414 -10 415 -9
rect 415 -10 416 -9
rect 416 -10 417 -9
rect 417 -10 418 -9
rect 418 -10 419 -9
rect 419 -10 420 -9
rect 420 -10 421 -9
rect 421 -10 422 -9
rect 422 -10 423 -9
rect 423 -10 424 -9
rect 424 -10 425 -9
rect 425 -10 426 -9
rect 426 -10 427 -9
rect 427 -10 428 -9
rect 428 -10 429 -9
rect 429 -10 430 -9
rect 430 -10 431 -9
rect 431 -10 432 -9
rect 432 -10 433 -9
rect 433 -10 434 -9
rect 434 -10 435 -9
rect 435 -10 436 -9
rect 436 -10 437 -9
rect 437 -10 438 -9
rect 438 -10 439 -9
rect 439 -10 440 -9
rect 440 -10 441 -9
rect 441 -10 442 -9
rect 442 -10 443 -9
rect 443 -10 444 -9
rect 444 -10 445 -9
rect 445 -10 446 -9
rect 446 -10 447 -9
rect 447 -10 448 -9
rect 448 -10 449 -9
rect 449 -10 450 -9
rect 450 -10 451 -9
rect 451 -10 452 -9
rect 452 -10 453 -9
rect 453 -10 454 -9
rect 454 -10 455 -9
rect 455 -10 456 -9
rect 456 -10 457 -9
rect 457 -10 458 -9
rect 458 -10 459 -9
rect 459 -10 460 -9
rect 460 -10 461 -9
rect 461 -10 462 -9
rect 462 -10 463 -9
rect 463 -10 464 -9
rect 464 -10 465 -9
rect 465 -10 466 -9
rect 466 -10 467 -9
rect 467 -10 468 -9
rect 468 -10 469 -9
rect 469 -10 470 -9
rect 470 -10 471 -9
rect 471 -10 472 -9
rect 472 -10 473 -9
rect 473 -10 474 -9
rect 474 -10 475 -9
rect 475 -10 476 -9
rect 476 -10 477 -9
rect 477 -10 478 -9
rect 478 -10 479 -9
rect 479 -10 480 -9
rect 2 -11 3 -10
rect 3 -11 4 -10
rect 4 -11 5 -10
rect 5 -11 6 -10
rect 6 -11 7 -10
rect 7 -11 8 -10
rect 8 -11 9 -10
rect 25 -11 26 -10
rect 26 -11 27 -10
rect 27 -11 28 -10
rect 28 -11 29 -10
rect 29 -11 30 -10
rect 30 -11 31 -10
rect 31 -11 32 -10
rect 32 -11 33 -10
rect 33 -11 34 -10
rect 34 -11 35 -10
rect 35 -11 36 -10
rect 36 -11 37 -10
rect 37 -11 38 -10
rect 38 -11 39 -10
rect 39 -11 40 -10
rect 40 -11 41 -10
rect 57 -11 58 -10
rect 58 -11 59 -10
rect 59 -11 60 -10
rect 60 -11 61 -10
rect 61 -11 62 -10
rect 62 -11 63 -10
rect 63 -11 64 -10
rect 64 -11 65 -10
rect 65 -11 66 -10
rect 66 -11 67 -10
rect 67 -11 68 -10
rect 68 -11 69 -10
rect 69 -11 70 -10
rect 70 -11 71 -10
rect 71 -11 72 -10
rect 72 -11 73 -10
rect 89 -11 90 -10
rect 90 -11 91 -10
rect 91 -11 92 -10
rect 92 -11 93 -10
rect 93 -11 94 -10
rect 94 -11 95 -10
rect 95 -11 96 -10
rect 96 -11 97 -10
rect 97 -11 98 -10
rect 98 -11 99 -10
rect 99 -11 100 -10
rect 100 -11 101 -10
rect 101 -11 102 -10
rect 102 -11 103 -10
rect 103 -11 104 -10
rect 104 -11 105 -10
rect 121 -11 122 -10
rect 122 -11 123 -10
rect 123 -11 124 -10
rect 124 -11 125 -10
rect 125 -11 126 -10
rect 126 -11 127 -10
rect 127 -11 128 -10
rect 128 -11 129 -10
rect 129 -11 130 -10
rect 130 -11 131 -10
rect 131 -11 132 -10
rect 132 -11 133 -10
rect 133 -11 134 -10
rect 134 -11 135 -10
rect 135 -11 136 -10
rect 136 -11 137 -10
rect 153 -11 154 -10
rect 154 -11 155 -10
rect 155 -11 156 -10
rect 156 -11 157 -10
rect 157 -11 158 -10
rect 158 -11 159 -10
rect 159 -11 160 -10
rect 160 -11 161 -10
rect 161 -11 162 -10
rect 162 -11 163 -10
rect 163 -11 164 -10
rect 164 -11 165 -10
rect 165 -11 166 -10
rect 166 -11 167 -10
rect 167 -11 168 -10
rect 168 -11 169 -10
rect 185 -11 186 -10
rect 186 -11 187 -10
rect 187 -11 188 -10
rect 188 -11 189 -10
rect 189 -11 190 -10
rect 190 -11 191 -10
rect 191 -11 192 -10
rect 192 -11 193 -10
rect 193 -11 194 -10
rect 194 -11 195 -10
rect 195 -11 196 -10
rect 196 -11 197 -10
rect 197 -11 198 -10
rect 198 -11 199 -10
rect 199 -11 200 -10
rect 200 -11 201 -10
rect 201 -11 202 -10
rect 202 -11 203 -10
rect 203 -11 204 -10
rect 204 -11 205 -10
rect 205 -11 206 -10
rect 206 -11 207 -10
rect 207 -11 208 -10
rect 208 -11 209 -10
rect 209 -11 210 -10
rect 210 -11 211 -10
rect 211 -11 212 -10
rect 212 -11 213 -10
rect 213 -11 214 -10
rect 214 -11 215 -10
rect 215 -11 216 -10
rect 216 -11 217 -10
rect 217 -11 218 -10
rect 218 -11 219 -10
rect 219 -11 220 -10
rect 220 -11 221 -10
rect 221 -11 222 -10
rect 222 -11 223 -10
rect 223 -11 224 -10
rect 224 -11 225 -10
rect 225 -11 226 -10
rect 226 -11 227 -10
rect 227 -11 228 -10
rect 228 -11 229 -10
rect 229 -11 230 -10
rect 230 -11 231 -10
rect 231 -11 232 -10
rect 232 -11 233 -10
rect 233 -11 234 -10
rect 234 -11 235 -10
rect 235 -11 236 -10
rect 236 -11 237 -10
rect 237 -11 238 -10
rect 238 -11 239 -10
rect 239 -11 240 -10
rect 240 -11 241 -10
rect 241 -11 242 -10
rect 242 -11 243 -10
rect 243 -11 244 -10
rect 244 -11 245 -10
rect 245 -11 246 -10
rect 246 -11 247 -10
rect 247 -11 248 -10
rect 248 -11 249 -10
rect 249 -11 250 -10
rect 250 -11 251 -10
rect 251 -11 252 -10
rect 252 -11 253 -10
rect 253 -11 254 -10
rect 254 -11 255 -10
rect 255 -11 256 -10
rect 256 -11 257 -10
rect 257 -11 258 -10
rect 258 -11 259 -10
rect 259 -11 260 -10
rect 260 -11 261 -10
rect 261 -11 262 -10
rect 262 -11 263 -10
rect 263 -11 264 -10
rect 264 -11 265 -10
rect 265 -11 266 -10
rect 266 -11 267 -10
rect 267 -11 268 -10
rect 268 -11 269 -10
rect 269 -11 270 -10
rect 270 -11 271 -10
rect 271 -11 272 -10
rect 272 -11 273 -10
rect 273 -11 274 -10
rect 274 -11 275 -10
rect 275 -11 276 -10
rect 276 -11 277 -10
rect 277 -11 278 -10
rect 278 -11 279 -10
rect 279 -11 280 -10
rect 280 -11 281 -10
rect 281 -11 282 -10
rect 282 -11 283 -10
rect 283 -11 284 -10
rect 284 -11 285 -10
rect 285 -11 286 -10
rect 286 -11 287 -10
rect 287 -11 288 -10
rect 288 -11 289 -10
rect 289 -11 290 -10
rect 290 -11 291 -10
rect 291 -11 292 -10
rect 292 -11 293 -10
rect 293 -11 294 -10
rect 294 -11 295 -10
rect 295 -11 296 -10
rect 296 -11 297 -10
rect 297 -11 298 -10
rect 298 -11 299 -10
rect 299 -11 300 -10
rect 300 -11 301 -10
rect 301 -11 302 -10
rect 302 -11 303 -10
rect 303 -11 304 -10
rect 304 -11 305 -10
rect 305 -11 306 -10
rect 306 -11 307 -10
rect 307 -11 308 -10
rect 308 -11 309 -10
rect 309 -11 310 -10
rect 310 -11 311 -10
rect 311 -11 312 -10
rect 312 -11 313 -10
rect 313 -11 314 -10
rect 314 -11 315 -10
rect 315 -11 316 -10
rect 316 -11 317 -10
rect 317 -11 318 -10
rect 318 -11 319 -10
rect 319 -11 320 -10
rect 320 -11 321 -10
rect 321 -11 322 -10
rect 322 -11 323 -10
rect 323 -11 324 -10
rect 324 -11 325 -10
rect 325 -11 326 -10
rect 326 -11 327 -10
rect 327 -11 328 -10
rect 328 -11 329 -10
rect 329 -11 330 -10
rect 330 -11 331 -10
rect 331 -11 332 -10
rect 332 -11 333 -10
rect 333 -11 334 -10
rect 334 -11 335 -10
rect 335 -11 336 -10
rect 336 -11 337 -10
rect 337 -11 338 -10
rect 338 -11 339 -10
rect 339 -11 340 -10
rect 340 -11 341 -10
rect 341 -11 342 -10
rect 342 -11 343 -10
rect 343 -11 344 -10
rect 344 -11 345 -10
rect 345 -11 346 -10
rect 346 -11 347 -10
rect 347 -11 348 -10
rect 348 -11 349 -10
rect 349 -11 350 -10
rect 350 -11 351 -10
rect 351 -11 352 -10
rect 352 -11 353 -10
rect 353 -11 354 -10
rect 354 -11 355 -10
rect 355 -11 356 -10
rect 356 -11 357 -10
rect 357 -11 358 -10
rect 358 -11 359 -10
rect 359 -11 360 -10
rect 360 -11 361 -10
rect 361 -11 362 -10
rect 362 -11 363 -10
rect 363 -11 364 -10
rect 364 -11 365 -10
rect 365 -11 366 -10
rect 366 -11 367 -10
rect 367 -11 368 -10
rect 368 -11 369 -10
rect 369 -11 370 -10
rect 370 -11 371 -10
rect 371 -11 372 -10
rect 372 -11 373 -10
rect 373 -11 374 -10
rect 374 -11 375 -10
rect 375 -11 376 -10
rect 376 -11 377 -10
rect 377 -11 378 -10
rect 378 -11 379 -10
rect 379 -11 380 -10
rect 380 -11 381 -10
rect 381 -11 382 -10
rect 382 -11 383 -10
rect 383 -11 384 -10
rect 384 -11 385 -10
rect 385 -11 386 -10
rect 386 -11 387 -10
rect 387 -11 388 -10
rect 388 -11 389 -10
rect 389 -11 390 -10
rect 390 -11 391 -10
rect 391 -11 392 -10
rect 392 -11 393 -10
rect 393 -11 394 -10
rect 394 -11 395 -10
rect 395 -11 396 -10
rect 396 -11 397 -10
rect 397 -11 398 -10
rect 398 -11 399 -10
rect 399 -11 400 -10
rect 400 -11 401 -10
rect 401 -11 402 -10
rect 402 -11 403 -10
rect 403 -11 404 -10
rect 404 -11 405 -10
rect 405 -11 406 -10
rect 406 -11 407 -10
rect 407 -11 408 -10
rect 408 -11 409 -10
rect 409 -11 410 -10
rect 410 -11 411 -10
rect 411 -11 412 -10
rect 412 -11 413 -10
rect 413 -11 414 -10
rect 414 -11 415 -10
rect 415 -11 416 -10
rect 416 -11 417 -10
rect 417 -11 418 -10
rect 418 -11 419 -10
rect 419 -11 420 -10
rect 420 -11 421 -10
rect 421 -11 422 -10
rect 422 -11 423 -10
rect 423 -11 424 -10
rect 424 -11 425 -10
rect 425 -11 426 -10
rect 426 -11 427 -10
rect 427 -11 428 -10
rect 428 -11 429 -10
rect 429 -11 430 -10
rect 430 -11 431 -10
rect 431 -11 432 -10
rect 432 -11 433 -10
rect 433 -11 434 -10
rect 434 -11 435 -10
rect 435 -11 436 -10
rect 436 -11 437 -10
rect 437 -11 438 -10
rect 438 -11 439 -10
rect 439 -11 440 -10
rect 440 -11 441 -10
rect 441 -11 442 -10
rect 442 -11 443 -10
rect 443 -11 444 -10
rect 444 -11 445 -10
rect 445 -11 446 -10
rect 446 -11 447 -10
rect 447 -11 448 -10
rect 448 -11 449 -10
rect 449 -11 450 -10
rect 450 -11 451 -10
rect 451 -11 452 -10
rect 452 -11 453 -10
rect 453 -11 454 -10
rect 454 -11 455 -10
rect 455 -11 456 -10
rect 456 -11 457 -10
rect 457 -11 458 -10
rect 458 -11 459 -10
rect 459 -11 460 -10
rect 460 -11 461 -10
rect 461 -11 462 -10
rect 462 -11 463 -10
rect 463 -11 464 -10
rect 464 -11 465 -10
rect 465 -11 466 -10
rect 466 -11 467 -10
rect 467 -11 468 -10
rect 468 -11 469 -10
rect 469 -11 470 -10
rect 470 -11 471 -10
rect 471 -11 472 -10
rect 472 -11 473 -10
rect 473 -11 474 -10
rect 474 -11 475 -10
rect 475 -11 476 -10
rect 476 -11 477 -10
rect 477 -11 478 -10
rect 478 -11 479 -10
rect 479 -11 480 -10
rect 2 -12 3 -11
rect 3 -12 4 -11
rect 4 -12 5 -11
rect 5 -12 6 -11
rect 6 -12 7 -11
rect 7 -12 8 -11
rect 8 -12 9 -11
rect 24 -12 25 -11
rect 25 -12 26 -11
rect 26 -12 27 -11
rect 27 -12 28 -11
rect 28 -12 29 -11
rect 29 -12 30 -11
rect 30 -12 31 -11
rect 31 -12 32 -11
rect 32 -12 33 -11
rect 33 -12 34 -11
rect 34 -12 35 -11
rect 35 -12 36 -11
rect 36 -12 37 -11
rect 37 -12 38 -11
rect 38 -12 39 -11
rect 39 -12 40 -11
rect 40 -12 41 -11
rect 56 -12 57 -11
rect 57 -12 58 -11
rect 58 -12 59 -11
rect 59 -12 60 -11
rect 60 -12 61 -11
rect 61 -12 62 -11
rect 62 -12 63 -11
rect 63 -12 64 -11
rect 64 -12 65 -11
rect 65 -12 66 -11
rect 66 -12 67 -11
rect 67 -12 68 -11
rect 68 -12 69 -11
rect 69 -12 70 -11
rect 70 -12 71 -11
rect 71 -12 72 -11
rect 72 -12 73 -11
rect 88 -12 89 -11
rect 89 -12 90 -11
rect 90 -12 91 -11
rect 91 -12 92 -11
rect 92 -12 93 -11
rect 93 -12 94 -11
rect 94 -12 95 -11
rect 95 -12 96 -11
rect 96 -12 97 -11
rect 97 -12 98 -11
rect 98 -12 99 -11
rect 99 -12 100 -11
rect 100 -12 101 -11
rect 101 -12 102 -11
rect 102 -12 103 -11
rect 103 -12 104 -11
rect 104 -12 105 -11
rect 120 -12 121 -11
rect 121 -12 122 -11
rect 122 -12 123 -11
rect 123 -12 124 -11
rect 124 -12 125 -11
rect 125 -12 126 -11
rect 126 -12 127 -11
rect 127 -12 128 -11
rect 128 -12 129 -11
rect 129 -12 130 -11
rect 130 -12 131 -11
rect 131 -12 132 -11
rect 132 -12 133 -11
rect 133 -12 134 -11
rect 134 -12 135 -11
rect 135 -12 136 -11
rect 136 -12 137 -11
rect 152 -12 153 -11
rect 153 -12 154 -11
rect 154 -12 155 -11
rect 155 -12 156 -11
rect 156 -12 157 -11
rect 157 -12 158 -11
rect 158 -12 159 -11
rect 159 -12 160 -11
rect 160 -12 161 -11
rect 161 -12 162 -11
rect 162 -12 163 -11
rect 163 -12 164 -11
rect 164 -12 165 -11
rect 165 -12 166 -11
rect 166 -12 167 -11
rect 167 -12 168 -11
rect 168 -12 169 -11
rect 184 -12 185 -11
rect 185 -12 186 -11
rect 186 -12 187 -11
rect 187 -12 188 -11
rect 188 -12 189 -11
rect 189 -12 190 -11
rect 190 -12 191 -11
rect 191 -12 192 -11
rect 192 -12 193 -11
rect 193 -12 194 -11
rect 194 -12 195 -11
rect 195 -12 196 -11
rect 196 -12 197 -11
rect 197 -12 198 -11
rect 198 -12 199 -11
rect 199 -12 200 -11
rect 200 -12 201 -11
rect 201 -12 202 -11
rect 202 -12 203 -11
rect 203 -12 204 -11
rect 204 -12 205 -11
rect 205 -12 206 -11
rect 206 -12 207 -11
rect 207 -12 208 -11
rect 208 -12 209 -11
rect 209 -12 210 -11
rect 210 -12 211 -11
rect 211 -12 212 -11
rect 212 -12 213 -11
rect 213 -12 214 -11
rect 214 -12 215 -11
rect 215 -12 216 -11
rect 216 -12 217 -11
rect 217 -12 218 -11
rect 218 -12 219 -11
rect 219 -12 220 -11
rect 220 -12 221 -11
rect 221 -12 222 -11
rect 222 -12 223 -11
rect 223 -12 224 -11
rect 224 -12 225 -11
rect 225 -12 226 -11
rect 226 -12 227 -11
rect 227 -12 228 -11
rect 228 -12 229 -11
rect 229 -12 230 -11
rect 230 -12 231 -11
rect 231 -12 232 -11
rect 232 -12 233 -11
rect 233 -12 234 -11
rect 234 -12 235 -11
rect 235 -12 236 -11
rect 236 -12 237 -11
rect 237 -12 238 -11
rect 238 -12 239 -11
rect 239 -12 240 -11
rect 240 -12 241 -11
rect 241 -12 242 -11
rect 242 -12 243 -11
rect 243 -12 244 -11
rect 244 -12 245 -11
rect 245 -12 246 -11
rect 246 -12 247 -11
rect 247 -12 248 -11
rect 248 -12 249 -11
rect 249 -12 250 -11
rect 250 -12 251 -11
rect 251 -12 252 -11
rect 252 -12 253 -11
rect 253 -12 254 -11
rect 254 -12 255 -11
rect 255 -12 256 -11
rect 256 -12 257 -11
rect 257 -12 258 -11
rect 258 -12 259 -11
rect 259 -12 260 -11
rect 260 -12 261 -11
rect 261 -12 262 -11
rect 262 -12 263 -11
rect 263 -12 264 -11
rect 264 -12 265 -11
rect 265 -12 266 -11
rect 266 -12 267 -11
rect 267 -12 268 -11
rect 268 -12 269 -11
rect 269 -12 270 -11
rect 270 -12 271 -11
rect 271 -12 272 -11
rect 272 -12 273 -11
rect 273 -12 274 -11
rect 274 -12 275 -11
rect 275 -12 276 -11
rect 276 -12 277 -11
rect 277 -12 278 -11
rect 278 -12 279 -11
rect 279 -12 280 -11
rect 280 -12 281 -11
rect 281 -12 282 -11
rect 282 -12 283 -11
rect 283 -12 284 -11
rect 284 -12 285 -11
rect 285 -12 286 -11
rect 286 -12 287 -11
rect 287 -12 288 -11
rect 288 -12 289 -11
rect 289 -12 290 -11
rect 290 -12 291 -11
rect 291 -12 292 -11
rect 292 -12 293 -11
rect 293 -12 294 -11
rect 294 -12 295 -11
rect 295 -12 296 -11
rect 296 -12 297 -11
rect 297 -12 298 -11
rect 298 -12 299 -11
rect 299 -12 300 -11
rect 300 -12 301 -11
rect 301 -12 302 -11
rect 302 -12 303 -11
rect 303 -12 304 -11
rect 304 -12 305 -11
rect 305 -12 306 -11
rect 306 -12 307 -11
rect 307 -12 308 -11
rect 308 -12 309 -11
rect 309 -12 310 -11
rect 310 -12 311 -11
rect 311 -12 312 -11
rect 312 -12 313 -11
rect 313 -12 314 -11
rect 314 -12 315 -11
rect 315 -12 316 -11
rect 316 -12 317 -11
rect 317 -12 318 -11
rect 318 -12 319 -11
rect 319 -12 320 -11
rect 320 -12 321 -11
rect 321 -12 322 -11
rect 322 -12 323 -11
rect 323 -12 324 -11
rect 324 -12 325 -11
rect 325 -12 326 -11
rect 326 -12 327 -11
rect 327 -12 328 -11
rect 328 -12 329 -11
rect 329 -12 330 -11
rect 330 -12 331 -11
rect 331 -12 332 -11
rect 332 -12 333 -11
rect 333 -12 334 -11
rect 334 -12 335 -11
rect 335 -12 336 -11
rect 336 -12 337 -11
rect 337 -12 338 -11
rect 338 -12 339 -11
rect 339 -12 340 -11
rect 340 -12 341 -11
rect 341 -12 342 -11
rect 342 -12 343 -11
rect 343 -12 344 -11
rect 344 -12 345 -11
rect 345 -12 346 -11
rect 346 -12 347 -11
rect 347 -12 348 -11
rect 348 -12 349 -11
rect 349 -12 350 -11
rect 350 -12 351 -11
rect 351 -12 352 -11
rect 352 -12 353 -11
rect 353 -12 354 -11
rect 354 -12 355 -11
rect 355 -12 356 -11
rect 356 -12 357 -11
rect 357 -12 358 -11
rect 358 -12 359 -11
rect 359 -12 360 -11
rect 360 -12 361 -11
rect 361 -12 362 -11
rect 362 -12 363 -11
rect 363 -12 364 -11
rect 364 -12 365 -11
rect 365 -12 366 -11
rect 366 -12 367 -11
rect 367 -12 368 -11
rect 368 -12 369 -11
rect 369 -12 370 -11
rect 370 -12 371 -11
rect 371 -12 372 -11
rect 372 -12 373 -11
rect 373 -12 374 -11
rect 374 -12 375 -11
rect 375 -12 376 -11
rect 376 -12 377 -11
rect 377 -12 378 -11
rect 378 -12 379 -11
rect 379 -12 380 -11
rect 380 -12 381 -11
rect 381 -12 382 -11
rect 382 -12 383 -11
rect 383 -12 384 -11
rect 384 -12 385 -11
rect 385 -12 386 -11
rect 386 -12 387 -11
rect 387 -12 388 -11
rect 388 -12 389 -11
rect 389 -12 390 -11
rect 390 -12 391 -11
rect 391 -12 392 -11
rect 392 -12 393 -11
rect 393 -12 394 -11
rect 394 -12 395 -11
rect 395 -12 396 -11
rect 396 -12 397 -11
rect 397 -12 398 -11
rect 398 -12 399 -11
rect 399 -12 400 -11
rect 400 -12 401 -11
rect 401 -12 402 -11
rect 402 -12 403 -11
rect 403 -12 404 -11
rect 404 -12 405 -11
rect 405 -12 406 -11
rect 406 -12 407 -11
rect 407 -12 408 -11
rect 408 -12 409 -11
rect 409 -12 410 -11
rect 410 -12 411 -11
rect 411 -12 412 -11
rect 412 -12 413 -11
rect 413 -12 414 -11
rect 414 -12 415 -11
rect 415 -12 416 -11
rect 416 -12 417 -11
rect 417 -12 418 -11
rect 418 -12 419 -11
rect 419 -12 420 -11
rect 420 -12 421 -11
rect 421 -12 422 -11
rect 422 -12 423 -11
rect 423 -12 424 -11
rect 424 -12 425 -11
rect 425 -12 426 -11
rect 426 -12 427 -11
rect 427 -12 428 -11
rect 428 -12 429 -11
rect 429 -12 430 -11
rect 430 -12 431 -11
rect 431 -12 432 -11
rect 432 -12 433 -11
rect 433 -12 434 -11
rect 434 -12 435 -11
rect 435 -12 436 -11
rect 436 -12 437 -11
rect 437 -12 438 -11
rect 438 -12 439 -11
rect 439 -12 440 -11
rect 440 -12 441 -11
rect 441 -12 442 -11
rect 442 -12 443 -11
rect 443 -12 444 -11
rect 444 -12 445 -11
rect 445 -12 446 -11
rect 446 -12 447 -11
rect 447 -12 448 -11
rect 448 -12 449 -11
rect 449 -12 450 -11
rect 450 -12 451 -11
rect 451 -12 452 -11
rect 452 -12 453 -11
rect 453 -12 454 -11
rect 454 -12 455 -11
rect 455 -12 456 -11
rect 456 -12 457 -11
rect 457 -12 458 -11
rect 458 -12 459 -11
rect 459 -12 460 -11
rect 460 -12 461 -11
rect 461 -12 462 -11
rect 462 -12 463 -11
rect 463 -12 464 -11
rect 464 -12 465 -11
rect 465 -12 466 -11
rect 466 -12 467 -11
rect 467 -12 468 -11
rect 468 -12 469 -11
rect 469 -12 470 -11
rect 470 -12 471 -11
rect 471 -12 472 -11
rect 472 -12 473 -11
rect 473 -12 474 -11
rect 474 -12 475 -11
rect 475 -12 476 -11
rect 476 -12 477 -11
rect 477 -12 478 -11
rect 478 -12 479 -11
rect 479 -12 480 -11
rect 2 -13 3 -12
rect 3 -13 4 -12
rect 4 -13 5 -12
rect 5 -13 6 -12
rect 6 -13 7 -12
rect 7 -13 8 -12
rect 8 -13 9 -12
rect 9 -13 10 -12
rect 10 -13 11 -12
rect 23 -13 24 -12
rect 24 -13 25 -12
rect 25 -13 26 -12
rect 26 -13 27 -12
rect 27 -13 28 -12
rect 28 -13 29 -12
rect 29 -13 30 -12
rect 30 -13 31 -12
rect 31 -13 32 -12
rect 32 -13 33 -12
rect 33 -13 34 -12
rect 34 -13 35 -12
rect 35 -13 36 -12
rect 36 -13 37 -12
rect 37 -13 38 -12
rect 38 -13 39 -12
rect 39 -13 40 -12
rect 40 -13 41 -12
rect 41 -13 42 -12
rect 42 -13 43 -12
rect 55 -13 56 -12
rect 56 -13 57 -12
rect 57 -13 58 -12
rect 58 -13 59 -12
rect 59 -13 60 -12
rect 60 -13 61 -12
rect 61 -13 62 -12
rect 62 -13 63 -12
rect 63 -13 64 -12
rect 64 -13 65 -12
rect 65 -13 66 -12
rect 66 -13 67 -12
rect 67 -13 68 -12
rect 68 -13 69 -12
rect 69 -13 70 -12
rect 70 -13 71 -12
rect 71 -13 72 -12
rect 72 -13 73 -12
rect 73 -13 74 -12
rect 74 -13 75 -12
rect 87 -13 88 -12
rect 88 -13 89 -12
rect 89 -13 90 -12
rect 90 -13 91 -12
rect 91 -13 92 -12
rect 92 -13 93 -12
rect 93 -13 94 -12
rect 94 -13 95 -12
rect 95 -13 96 -12
rect 96 -13 97 -12
rect 97 -13 98 -12
rect 98 -13 99 -12
rect 99 -13 100 -12
rect 100 -13 101 -12
rect 101 -13 102 -12
rect 102 -13 103 -12
rect 103 -13 104 -12
rect 104 -13 105 -12
rect 105 -13 106 -12
rect 106 -13 107 -12
rect 119 -13 120 -12
rect 120 -13 121 -12
rect 121 -13 122 -12
rect 122 -13 123 -12
rect 123 -13 124 -12
rect 124 -13 125 -12
rect 125 -13 126 -12
rect 126 -13 127 -12
rect 127 -13 128 -12
rect 128 -13 129 -12
rect 129 -13 130 -12
rect 130 -13 131 -12
rect 131 -13 132 -12
rect 132 -13 133 -12
rect 133 -13 134 -12
rect 134 -13 135 -12
rect 135 -13 136 -12
rect 136 -13 137 -12
rect 137 -13 138 -12
rect 138 -13 139 -12
rect 151 -13 152 -12
rect 152 -13 153 -12
rect 153 -13 154 -12
rect 154 -13 155 -12
rect 155 -13 156 -12
rect 156 -13 157 -12
rect 157 -13 158 -12
rect 158 -13 159 -12
rect 159 -13 160 -12
rect 160 -13 161 -12
rect 161 -13 162 -12
rect 162 -13 163 -12
rect 163 -13 164 -12
rect 164 -13 165 -12
rect 165 -13 166 -12
rect 166 -13 167 -12
rect 167 -13 168 -12
rect 168 -13 169 -12
rect 169 -13 170 -12
rect 170 -13 171 -12
rect 183 -13 184 -12
rect 184 -13 185 -12
rect 185 -13 186 -12
rect 186 -13 187 -12
rect 187 -13 188 -12
rect 188 -13 189 -12
rect 189 -13 190 -12
rect 190 -13 191 -12
rect 191 -13 192 -12
rect 192 -13 193 -12
rect 193 -13 194 -12
rect 194 -13 195 -12
rect 195 -13 196 -12
rect 196 -13 197 -12
rect 197 -13 198 -12
rect 198 -13 199 -12
rect 199 -13 200 -12
rect 200 -13 201 -12
rect 201 -13 202 -12
rect 202 -13 203 -12
rect 203 -13 204 -12
rect 204 -13 205 -12
rect 205 -13 206 -12
rect 206 -13 207 -12
rect 207 -13 208 -12
rect 208 -13 209 -12
rect 209 -13 210 -12
rect 210 -13 211 -12
rect 211 -13 212 -12
rect 212 -13 213 -12
rect 213 -13 214 -12
rect 214 -13 215 -12
rect 215 -13 216 -12
rect 216 -13 217 -12
rect 217 -13 218 -12
rect 218 -13 219 -12
rect 219 -13 220 -12
rect 220 -13 221 -12
rect 221 -13 222 -12
rect 222 -13 223 -12
rect 223 -13 224 -12
rect 224 -13 225 -12
rect 225 -13 226 -12
rect 226 -13 227 -12
rect 227 -13 228 -12
rect 228 -13 229 -12
rect 229 -13 230 -12
rect 230 -13 231 -12
rect 231 -13 232 -12
rect 232 -13 233 -12
rect 233 -13 234 -12
rect 234 -13 235 -12
rect 235 -13 236 -12
rect 236 -13 237 -12
rect 237 -13 238 -12
rect 238 -13 239 -12
rect 239 -13 240 -12
rect 240 -13 241 -12
rect 241 -13 242 -12
rect 242 -13 243 -12
rect 243 -13 244 -12
rect 244 -13 245 -12
rect 245 -13 246 -12
rect 246 -13 247 -12
rect 247 -13 248 -12
rect 248 -13 249 -12
rect 249 -13 250 -12
rect 250 -13 251 -12
rect 251 -13 252 -12
rect 252 -13 253 -12
rect 253 -13 254 -12
rect 254 -13 255 -12
rect 255 -13 256 -12
rect 256 -13 257 -12
rect 257 -13 258 -12
rect 258 -13 259 -12
rect 259 -13 260 -12
rect 260 -13 261 -12
rect 261 -13 262 -12
rect 262 -13 263 -12
rect 263 -13 264 -12
rect 264 -13 265 -12
rect 265 -13 266 -12
rect 266 -13 267 -12
rect 267 -13 268 -12
rect 268 -13 269 -12
rect 269 -13 270 -12
rect 270 -13 271 -12
rect 271 -13 272 -12
rect 272 -13 273 -12
rect 273 -13 274 -12
rect 274 -13 275 -12
rect 275 -13 276 -12
rect 276 -13 277 -12
rect 277 -13 278 -12
rect 278 -13 279 -12
rect 279 -13 280 -12
rect 280 -13 281 -12
rect 281 -13 282 -12
rect 282 -13 283 -12
rect 283 -13 284 -12
rect 284 -13 285 -12
rect 285 -13 286 -12
rect 286 -13 287 -12
rect 287 -13 288 -12
rect 288 -13 289 -12
rect 289 -13 290 -12
rect 290 -13 291 -12
rect 291 -13 292 -12
rect 292 -13 293 -12
rect 293 -13 294 -12
rect 294 -13 295 -12
rect 295 -13 296 -12
rect 296 -13 297 -12
rect 297 -13 298 -12
rect 298 -13 299 -12
rect 299 -13 300 -12
rect 300 -13 301 -12
rect 301 -13 302 -12
rect 302 -13 303 -12
rect 303 -13 304 -12
rect 304 -13 305 -12
rect 305 -13 306 -12
rect 306 -13 307 -12
rect 307 -13 308 -12
rect 308 -13 309 -12
rect 309 -13 310 -12
rect 310 -13 311 -12
rect 311 -13 312 -12
rect 312 -13 313 -12
rect 313 -13 314 -12
rect 314 -13 315 -12
rect 315 -13 316 -12
rect 316 -13 317 -12
rect 317 -13 318 -12
rect 318 -13 319 -12
rect 319 -13 320 -12
rect 320 -13 321 -12
rect 321 -13 322 -12
rect 322 -13 323 -12
rect 323 -13 324 -12
rect 324 -13 325 -12
rect 325 -13 326 -12
rect 326 -13 327 -12
rect 327 -13 328 -12
rect 328 -13 329 -12
rect 329 -13 330 -12
rect 330 -13 331 -12
rect 331 -13 332 -12
rect 332 -13 333 -12
rect 333 -13 334 -12
rect 334 -13 335 -12
rect 335 -13 336 -12
rect 336 -13 337 -12
rect 337 -13 338 -12
rect 338 -13 339 -12
rect 339 -13 340 -12
rect 340 -13 341 -12
rect 341 -13 342 -12
rect 342 -13 343 -12
rect 343 -13 344 -12
rect 344 -13 345 -12
rect 345 -13 346 -12
rect 346 -13 347 -12
rect 347 -13 348 -12
rect 348 -13 349 -12
rect 349 -13 350 -12
rect 350 -13 351 -12
rect 351 -13 352 -12
rect 352 -13 353 -12
rect 353 -13 354 -12
rect 354 -13 355 -12
rect 355 -13 356 -12
rect 356 -13 357 -12
rect 357 -13 358 -12
rect 358 -13 359 -12
rect 359 -13 360 -12
rect 360 -13 361 -12
rect 361 -13 362 -12
rect 362 -13 363 -12
rect 363 -13 364 -12
rect 364 -13 365 -12
rect 365 -13 366 -12
rect 366 -13 367 -12
rect 367 -13 368 -12
rect 368 -13 369 -12
rect 369 -13 370 -12
rect 370 -13 371 -12
rect 371 -13 372 -12
rect 372 -13 373 -12
rect 373 -13 374 -12
rect 374 -13 375 -12
rect 375 -13 376 -12
rect 376 -13 377 -12
rect 377 -13 378 -12
rect 378 -13 379 -12
rect 379 -13 380 -12
rect 380 -13 381 -12
rect 381 -13 382 -12
rect 382 -13 383 -12
rect 383 -13 384 -12
rect 384 -13 385 -12
rect 385 -13 386 -12
rect 386 -13 387 -12
rect 387 -13 388 -12
rect 388 -13 389 -12
rect 389 -13 390 -12
rect 390 -13 391 -12
rect 391 -13 392 -12
rect 392 -13 393 -12
rect 393 -13 394 -12
rect 394 -13 395 -12
rect 395 -13 396 -12
rect 396 -13 397 -12
rect 397 -13 398 -12
rect 398 -13 399 -12
rect 399 -13 400 -12
rect 400 -13 401 -12
rect 401 -13 402 -12
rect 402 -13 403 -12
rect 403 -13 404 -12
rect 404 -13 405 -12
rect 405 -13 406 -12
rect 406 -13 407 -12
rect 407 -13 408 -12
rect 408 -13 409 -12
rect 409 -13 410 -12
rect 410 -13 411 -12
rect 411 -13 412 -12
rect 412 -13 413 -12
rect 413 -13 414 -12
rect 414 -13 415 -12
rect 415 -13 416 -12
rect 416 -13 417 -12
rect 417 -13 418 -12
rect 418 -13 419 -12
rect 419 -13 420 -12
rect 420 -13 421 -12
rect 421 -13 422 -12
rect 422 -13 423 -12
rect 423 -13 424 -12
rect 424 -13 425 -12
rect 425 -13 426 -12
rect 426 -13 427 -12
rect 427 -13 428 -12
rect 428 -13 429 -12
rect 429 -13 430 -12
rect 430 -13 431 -12
rect 431 -13 432 -12
rect 432 -13 433 -12
rect 433 -13 434 -12
rect 434 -13 435 -12
rect 435 -13 436 -12
rect 436 -13 437 -12
rect 437 -13 438 -12
rect 438 -13 439 -12
rect 439 -13 440 -12
rect 440 -13 441 -12
rect 441 -13 442 -12
rect 442 -13 443 -12
rect 443 -13 444 -12
rect 444 -13 445 -12
rect 445 -13 446 -12
rect 446 -13 447 -12
rect 447 -13 448 -12
rect 448 -13 449 -12
rect 449 -13 450 -12
rect 450 -13 451 -12
rect 451 -13 452 -12
rect 452 -13 453 -12
rect 453 -13 454 -12
rect 454 -13 455 -12
rect 455 -13 456 -12
rect 456 -13 457 -12
rect 457 -13 458 -12
rect 458 -13 459 -12
rect 459 -13 460 -12
rect 460 -13 461 -12
rect 461 -13 462 -12
rect 462 -13 463 -12
rect 463 -13 464 -12
rect 464 -13 465 -12
rect 465 -13 466 -12
rect 466 -13 467 -12
rect 467 -13 468 -12
rect 468 -13 469 -12
rect 469 -13 470 -12
rect 470 -13 471 -12
rect 471 -13 472 -12
rect 472 -13 473 -12
rect 473 -13 474 -12
rect 474 -13 475 -12
rect 475 -13 476 -12
rect 476 -13 477 -12
rect 477 -13 478 -12
rect 478 -13 479 -12
rect 479 -13 480 -12
rect 2 -14 3 -13
rect 3 -14 4 -13
rect 4 -14 5 -13
rect 5 -14 6 -13
rect 6 -14 7 -13
rect 7 -14 8 -13
rect 8 -14 9 -13
rect 9 -14 10 -13
rect 10 -14 11 -13
rect 11 -14 12 -13
rect 22 -14 23 -13
rect 23 -14 24 -13
rect 24 -14 25 -13
rect 25 -14 26 -13
rect 26 -14 27 -13
rect 27 -14 28 -13
rect 28 -14 29 -13
rect 29 -14 30 -13
rect 30 -14 31 -13
rect 31 -14 32 -13
rect 32 -14 33 -13
rect 33 -14 34 -13
rect 34 -14 35 -13
rect 35 -14 36 -13
rect 36 -14 37 -13
rect 37 -14 38 -13
rect 38 -14 39 -13
rect 39 -14 40 -13
rect 40 -14 41 -13
rect 41 -14 42 -13
rect 42 -14 43 -13
rect 43 -14 44 -13
rect 54 -14 55 -13
rect 55 -14 56 -13
rect 56 -14 57 -13
rect 57 -14 58 -13
rect 58 -14 59 -13
rect 59 -14 60 -13
rect 60 -14 61 -13
rect 61 -14 62 -13
rect 62 -14 63 -13
rect 63 -14 64 -13
rect 64 -14 65 -13
rect 65 -14 66 -13
rect 66 -14 67 -13
rect 67 -14 68 -13
rect 68 -14 69 -13
rect 69 -14 70 -13
rect 70 -14 71 -13
rect 71 -14 72 -13
rect 72 -14 73 -13
rect 73 -14 74 -13
rect 74 -14 75 -13
rect 75 -14 76 -13
rect 86 -14 87 -13
rect 87 -14 88 -13
rect 88 -14 89 -13
rect 89 -14 90 -13
rect 90 -14 91 -13
rect 91 -14 92 -13
rect 92 -14 93 -13
rect 93 -14 94 -13
rect 94 -14 95 -13
rect 95 -14 96 -13
rect 96 -14 97 -13
rect 97 -14 98 -13
rect 98 -14 99 -13
rect 99 -14 100 -13
rect 100 -14 101 -13
rect 101 -14 102 -13
rect 102 -14 103 -13
rect 103 -14 104 -13
rect 104 -14 105 -13
rect 105 -14 106 -13
rect 106 -14 107 -13
rect 107 -14 108 -13
rect 118 -14 119 -13
rect 119 -14 120 -13
rect 120 -14 121 -13
rect 121 -14 122 -13
rect 122 -14 123 -13
rect 123 -14 124 -13
rect 124 -14 125 -13
rect 125 -14 126 -13
rect 126 -14 127 -13
rect 127 -14 128 -13
rect 128 -14 129 -13
rect 129 -14 130 -13
rect 130 -14 131 -13
rect 131 -14 132 -13
rect 132 -14 133 -13
rect 133 -14 134 -13
rect 134 -14 135 -13
rect 135 -14 136 -13
rect 136 -14 137 -13
rect 137 -14 138 -13
rect 138 -14 139 -13
rect 139 -14 140 -13
rect 150 -14 151 -13
rect 151 -14 152 -13
rect 152 -14 153 -13
rect 153 -14 154 -13
rect 154 -14 155 -13
rect 155 -14 156 -13
rect 156 -14 157 -13
rect 157 -14 158 -13
rect 158 -14 159 -13
rect 159 -14 160 -13
rect 160 -14 161 -13
rect 161 -14 162 -13
rect 162 -14 163 -13
rect 163 -14 164 -13
rect 164 -14 165 -13
rect 165 -14 166 -13
rect 166 -14 167 -13
rect 167 -14 168 -13
rect 168 -14 169 -13
rect 169 -14 170 -13
rect 170 -14 171 -13
rect 171 -14 172 -13
rect 182 -14 183 -13
rect 183 -14 184 -13
rect 184 -14 185 -13
rect 185 -14 186 -13
rect 186 -14 187 -13
rect 187 -14 188 -13
rect 188 -14 189 -13
rect 189 -14 190 -13
rect 190 -14 191 -13
rect 191 -14 192 -13
rect 192 -14 193 -13
rect 193 -14 194 -13
rect 194 -14 195 -13
rect 195 -14 196 -13
rect 196 -14 197 -13
rect 197 -14 198 -13
rect 198 -14 199 -13
rect 199 -14 200 -13
rect 200 -14 201 -13
rect 201 -14 202 -13
rect 202 -14 203 -13
rect 203 -14 204 -13
rect 204 -14 205 -13
rect 205 -14 206 -13
rect 206 -14 207 -13
rect 207 -14 208 -13
rect 208 -14 209 -13
rect 209 -14 210 -13
rect 210 -14 211 -13
rect 211 -14 212 -13
rect 212 -14 213 -13
rect 213 -14 214 -13
rect 214 -14 215 -13
rect 215 -14 216 -13
rect 216 -14 217 -13
rect 217 -14 218 -13
rect 218 -14 219 -13
rect 219 -14 220 -13
rect 220 -14 221 -13
rect 221 -14 222 -13
rect 222 -14 223 -13
rect 223 -14 224 -13
rect 224 -14 225 -13
rect 225 -14 226 -13
rect 226 -14 227 -13
rect 227 -14 228 -13
rect 228 -14 229 -13
rect 229 -14 230 -13
rect 230 -14 231 -13
rect 231 -14 232 -13
rect 232 -14 233 -13
rect 233 -14 234 -13
rect 234 -14 235 -13
rect 235 -14 236 -13
rect 236 -14 237 -13
rect 237 -14 238 -13
rect 238 -14 239 -13
rect 239 -14 240 -13
rect 240 -14 241 -13
rect 241 -14 242 -13
rect 242 -14 243 -13
rect 243 -14 244 -13
rect 244 -14 245 -13
rect 245 -14 246 -13
rect 246 -14 247 -13
rect 247 -14 248 -13
rect 248 -14 249 -13
rect 249 -14 250 -13
rect 250 -14 251 -13
rect 251 -14 252 -13
rect 252 -14 253 -13
rect 253 -14 254 -13
rect 254 -14 255 -13
rect 255 -14 256 -13
rect 256 -14 257 -13
rect 257 -14 258 -13
rect 258 -14 259 -13
rect 259 -14 260 -13
rect 260 -14 261 -13
rect 261 -14 262 -13
rect 262 -14 263 -13
rect 263 -14 264 -13
rect 264 -14 265 -13
rect 265 -14 266 -13
rect 266 -14 267 -13
rect 267 -14 268 -13
rect 268 -14 269 -13
rect 269 -14 270 -13
rect 270 -14 271 -13
rect 271 -14 272 -13
rect 272 -14 273 -13
rect 273 -14 274 -13
rect 274 -14 275 -13
rect 275 -14 276 -13
rect 276 -14 277 -13
rect 277 -14 278 -13
rect 278 -14 279 -13
rect 279 -14 280 -13
rect 280 -14 281 -13
rect 281 -14 282 -13
rect 282 -14 283 -13
rect 283 -14 284 -13
rect 284 -14 285 -13
rect 285 -14 286 -13
rect 286 -14 287 -13
rect 287 -14 288 -13
rect 288 -14 289 -13
rect 289 -14 290 -13
rect 290 -14 291 -13
rect 291 -14 292 -13
rect 292 -14 293 -13
rect 293 -14 294 -13
rect 294 -14 295 -13
rect 295 -14 296 -13
rect 296 -14 297 -13
rect 297 -14 298 -13
rect 298 -14 299 -13
rect 299 -14 300 -13
rect 300 -14 301 -13
rect 301 -14 302 -13
rect 302 -14 303 -13
rect 303 -14 304 -13
rect 304 -14 305 -13
rect 305 -14 306 -13
rect 306 -14 307 -13
rect 307 -14 308 -13
rect 308 -14 309 -13
rect 309 -14 310 -13
rect 310 -14 311 -13
rect 311 -14 312 -13
rect 312 -14 313 -13
rect 313 -14 314 -13
rect 314 -14 315 -13
rect 315 -14 316 -13
rect 316 -14 317 -13
rect 317 -14 318 -13
rect 318 -14 319 -13
rect 319 -14 320 -13
rect 320 -14 321 -13
rect 321 -14 322 -13
rect 322 -14 323 -13
rect 323 -14 324 -13
rect 324 -14 325 -13
rect 325 -14 326 -13
rect 326 -14 327 -13
rect 327 -14 328 -13
rect 328 -14 329 -13
rect 329 -14 330 -13
rect 330 -14 331 -13
rect 331 -14 332 -13
rect 332 -14 333 -13
rect 333 -14 334 -13
rect 334 -14 335 -13
rect 335 -14 336 -13
rect 336 -14 337 -13
rect 337 -14 338 -13
rect 338 -14 339 -13
rect 339 -14 340 -13
rect 340 -14 341 -13
rect 341 -14 342 -13
rect 342 -14 343 -13
rect 343 -14 344 -13
rect 344 -14 345 -13
rect 345 -14 346 -13
rect 346 -14 347 -13
rect 347 -14 348 -13
rect 348 -14 349 -13
rect 349 -14 350 -13
rect 350 -14 351 -13
rect 351 -14 352 -13
rect 352 -14 353 -13
rect 353 -14 354 -13
rect 354 -14 355 -13
rect 355 -14 356 -13
rect 356 -14 357 -13
rect 357 -14 358 -13
rect 358 -14 359 -13
rect 359 -14 360 -13
rect 360 -14 361 -13
rect 361 -14 362 -13
rect 362 -14 363 -13
rect 363 -14 364 -13
rect 364 -14 365 -13
rect 365 -14 366 -13
rect 366 -14 367 -13
rect 367 -14 368 -13
rect 368 -14 369 -13
rect 369 -14 370 -13
rect 370 -14 371 -13
rect 371 -14 372 -13
rect 372 -14 373 -13
rect 373 -14 374 -13
rect 374 -14 375 -13
rect 375 -14 376 -13
rect 376 -14 377 -13
rect 377 -14 378 -13
rect 378 -14 379 -13
rect 379 -14 380 -13
rect 380 -14 381 -13
rect 381 -14 382 -13
rect 382 -14 383 -13
rect 383 -14 384 -13
rect 384 -14 385 -13
rect 385 -14 386 -13
rect 386 -14 387 -13
rect 387 -14 388 -13
rect 388 -14 389 -13
rect 389 -14 390 -13
rect 390 -14 391 -13
rect 391 -14 392 -13
rect 392 -14 393 -13
rect 393 -14 394 -13
rect 394 -14 395 -13
rect 395 -14 396 -13
rect 396 -14 397 -13
rect 397 -14 398 -13
rect 398 -14 399 -13
rect 399 -14 400 -13
rect 400 -14 401 -13
rect 401 -14 402 -13
rect 402 -14 403 -13
rect 403 -14 404 -13
rect 404 -14 405 -13
rect 405 -14 406 -13
rect 406 -14 407 -13
rect 407 -14 408 -13
rect 408 -14 409 -13
rect 409 -14 410 -13
rect 410 -14 411 -13
rect 411 -14 412 -13
rect 412 -14 413 -13
rect 413 -14 414 -13
rect 414 -14 415 -13
rect 415 -14 416 -13
rect 416 -14 417 -13
rect 417 -14 418 -13
rect 418 -14 419 -13
rect 419 -14 420 -13
rect 420 -14 421 -13
rect 421 -14 422 -13
rect 422 -14 423 -13
rect 423 -14 424 -13
rect 424 -14 425 -13
rect 425 -14 426 -13
rect 426 -14 427 -13
rect 427 -14 428 -13
rect 428 -14 429 -13
rect 429 -14 430 -13
rect 430 -14 431 -13
rect 431 -14 432 -13
rect 432 -14 433 -13
rect 433 -14 434 -13
rect 434 -14 435 -13
rect 435 -14 436 -13
rect 436 -14 437 -13
rect 437 -14 438 -13
rect 438 -14 439 -13
rect 439 -14 440 -13
rect 440 -14 441 -13
rect 441 -14 442 -13
rect 442 -14 443 -13
rect 443 -14 444 -13
rect 444 -14 445 -13
rect 445 -14 446 -13
rect 446 -14 447 -13
rect 447 -14 448 -13
rect 448 -14 449 -13
rect 449 -14 450 -13
rect 450 -14 451 -13
rect 451 -14 452 -13
rect 452 -14 453 -13
rect 453 -14 454 -13
rect 454 -14 455 -13
rect 455 -14 456 -13
rect 456 -14 457 -13
rect 457 -14 458 -13
rect 458 -14 459 -13
rect 459 -14 460 -13
rect 460 -14 461 -13
rect 461 -14 462 -13
rect 462 -14 463 -13
rect 463 -14 464 -13
rect 464 -14 465 -13
rect 465 -14 466 -13
rect 466 -14 467 -13
rect 467 -14 468 -13
rect 468 -14 469 -13
rect 469 -14 470 -13
rect 470 -14 471 -13
rect 471 -14 472 -13
rect 472 -14 473 -13
rect 473 -14 474 -13
rect 474 -14 475 -13
rect 475 -14 476 -13
rect 476 -14 477 -13
rect 477 -14 478 -13
rect 478 -14 479 -13
rect 479 -14 480 -13
rect 2 -15 3 -14
rect 3 -15 4 -14
rect 4 -15 5 -14
rect 5 -15 6 -14
rect 6 -15 7 -14
rect 7 -15 8 -14
rect 8 -15 9 -14
rect 9 -15 10 -14
rect 10 -15 11 -14
rect 11 -15 12 -14
rect 21 -15 22 -14
rect 22 -15 23 -14
rect 23 -15 24 -14
rect 24 -15 25 -14
rect 25 -15 26 -14
rect 26 -15 27 -14
rect 27 -15 28 -14
rect 28 -15 29 -14
rect 29 -15 30 -14
rect 30 -15 31 -14
rect 31 -15 32 -14
rect 32 -15 33 -14
rect 33 -15 34 -14
rect 34 -15 35 -14
rect 35 -15 36 -14
rect 36 -15 37 -14
rect 37 -15 38 -14
rect 38 -15 39 -14
rect 39 -15 40 -14
rect 40 -15 41 -14
rect 41 -15 42 -14
rect 42 -15 43 -14
rect 43 -15 44 -14
rect 53 -15 54 -14
rect 54 -15 55 -14
rect 55 -15 56 -14
rect 56 -15 57 -14
rect 57 -15 58 -14
rect 58 -15 59 -14
rect 59 -15 60 -14
rect 60 -15 61 -14
rect 61 -15 62 -14
rect 62 -15 63 -14
rect 63 -15 64 -14
rect 64 -15 65 -14
rect 65 -15 66 -14
rect 66 -15 67 -14
rect 67 -15 68 -14
rect 68 -15 69 -14
rect 69 -15 70 -14
rect 70 -15 71 -14
rect 71 -15 72 -14
rect 72 -15 73 -14
rect 73 -15 74 -14
rect 74 -15 75 -14
rect 75 -15 76 -14
rect 85 -15 86 -14
rect 86 -15 87 -14
rect 87 -15 88 -14
rect 88 -15 89 -14
rect 89 -15 90 -14
rect 90 -15 91 -14
rect 91 -15 92 -14
rect 92 -15 93 -14
rect 93 -15 94 -14
rect 94 -15 95 -14
rect 95 -15 96 -14
rect 96 -15 97 -14
rect 97 -15 98 -14
rect 98 -15 99 -14
rect 99 -15 100 -14
rect 100 -15 101 -14
rect 101 -15 102 -14
rect 102 -15 103 -14
rect 103 -15 104 -14
rect 104 -15 105 -14
rect 105 -15 106 -14
rect 106 -15 107 -14
rect 107 -15 108 -14
rect 117 -15 118 -14
rect 118 -15 119 -14
rect 119 -15 120 -14
rect 120 -15 121 -14
rect 121 -15 122 -14
rect 122 -15 123 -14
rect 123 -15 124 -14
rect 124 -15 125 -14
rect 125 -15 126 -14
rect 126 -15 127 -14
rect 127 -15 128 -14
rect 128 -15 129 -14
rect 129 -15 130 -14
rect 130 -15 131 -14
rect 131 -15 132 -14
rect 132 -15 133 -14
rect 133 -15 134 -14
rect 134 -15 135 -14
rect 135 -15 136 -14
rect 136 -15 137 -14
rect 137 -15 138 -14
rect 138 -15 139 -14
rect 139 -15 140 -14
rect 149 -15 150 -14
rect 150 -15 151 -14
rect 151 -15 152 -14
rect 152 -15 153 -14
rect 153 -15 154 -14
rect 154 -15 155 -14
rect 155 -15 156 -14
rect 156 -15 157 -14
rect 157 -15 158 -14
rect 158 -15 159 -14
rect 159 -15 160 -14
rect 160 -15 161 -14
rect 161 -15 162 -14
rect 162 -15 163 -14
rect 163 -15 164 -14
rect 164 -15 165 -14
rect 165 -15 166 -14
rect 166 -15 167 -14
rect 167 -15 168 -14
rect 168 -15 169 -14
rect 169 -15 170 -14
rect 170 -15 171 -14
rect 171 -15 172 -14
rect 181 -15 182 -14
rect 182 -15 183 -14
rect 183 -15 184 -14
rect 184 -15 185 -14
rect 185 -15 186 -14
rect 186 -15 187 -14
rect 187 -15 188 -14
rect 188 -15 189 -14
rect 189 -15 190 -14
rect 190 -15 191 -14
rect 191 -15 192 -14
rect 192 -15 193 -14
rect 193 -15 194 -14
rect 194 -15 195 -14
rect 195 -15 196 -14
rect 196 -15 197 -14
rect 197 -15 198 -14
rect 198 -15 199 -14
rect 199 -15 200 -14
rect 200 -15 201 -14
rect 201 -15 202 -14
rect 202 -15 203 -14
rect 203 -15 204 -14
rect 204 -15 205 -14
rect 205 -15 206 -14
rect 206 -15 207 -14
rect 207 -15 208 -14
rect 208 -15 209 -14
rect 209 -15 210 -14
rect 210 -15 211 -14
rect 211 -15 212 -14
rect 212 -15 213 -14
rect 213 -15 214 -14
rect 214 -15 215 -14
rect 215 -15 216 -14
rect 216 -15 217 -14
rect 217 -15 218 -14
rect 218 -15 219 -14
rect 219 -15 220 -14
rect 220 -15 221 -14
rect 221 -15 222 -14
rect 222 -15 223 -14
rect 223 -15 224 -14
rect 224 -15 225 -14
rect 225 -15 226 -14
rect 226 -15 227 -14
rect 227 -15 228 -14
rect 228 -15 229 -14
rect 229 -15 230 -14
rect 230 -15 231 -14
rect 231 -15 232 -14
rect 232 -15 233 -14
rect 233 -15 234 -14
rect 234 -15 235 -14
rect 235 -15 236 -14
rect 236 -15 237 -14
rect 237 -15 238 -14
rect 238 -15 239 -14
rect 239 -15 240 -14
rect 240 -15 241 -14
rect 241 -15 242 -14
rect 242 -15 243 -14
rect 243 -15 244 -14
rect 244 -15 245 -14
rect 245 -15 246 -14
rect 246 -15 247 -14
rect 247 -15 248 -14
rect 248 -15 249 -14
rect 249 -15 250 -14
rect 250 -15 251 -14
rect 251 -15 252 -14
rect 252 -15 253 -14
rect 253 -15 254 -14
rect 254 -15 255 -14
rect 255 -15 256 -14
rect 256 -15 257 -14
rect 257 -15 258 -14
rect 258 -15 259 -14
rect 259 -15 260 -14
rect 260 -15 261 -14
rect 261 -15 262 -14
rect 262 -15 263 -14
rect 263 -15 264 -14
rect 264 -15 265 -14
rect 265 -15 266 -14
rect 266 -15 267 -14
rect 267 -15 268 -14
rect 268 -15 269 -14
rect 269 -15 270 -14
rect 270 -15 271 -14
rect 271 -15 272 -14
rect 272 -15 273 -14
rect 273 -15 274 -14
rect 274 -15 275 -14
rect 275 -15 276 -14
rect 276 -15 277 -14
rect 277 -15 278 -14
rect 278 -15 279 -14
rect 279 -15 280 -14
rect 280 -15 281 -14
rect 281 -15 282 -14
rect 282 -15 283 -14
rect 283 -15 284 -14
rect 284 -15 285 -14
rect 285 -15 286 -14
rect 286 -15 287 -14
rect 287 -15 288 -14
rect 288 -15 289 -14
rect 289 -15 290 -14
rect 290 -15 291 -14
rect 291 -15 292 -14
rect 292 -15 293 -14
rect 293 -15 294 -14
rect 294 -15 295 -14
rect 295 -15 296 -14
rect 296 -15 297 -14
rect 297 -15 298 -14
rect 298 -15 299 -14
rect 299 -15 300 -14
rect 300 -15 301 -14
rect 301 -15 302 -14
rect 302 -15 303 -14
rect 303 -15 304 -14
rect 304 -15 305 -14
rect 305 -15 306 -14
rect 306 -15 307 -14
rect 307 -15 308 -14
rect 308 -15 309 -14
rect 309 -15 310 -14
rect 310 -15 311 -14
rect 311 -15 312 -14
rect 312 -15 313 -14
rect 313 -15 314 -14
rect 314 -15 315 -14
rect 315 -15 316 -14
rect 316 -15 317 -14
rect 317 -15 318 -14
rect 318 -15 319 -14
rect 319 -15 320 -14
rect 320 -15 321 -14
rect 321 -15 322 -14
rect 322 -15 323 -14
rect 323 -15 324 -14
rect 324 -15 325 -14
rect 325 -15 326 -14
rect 326 -15 327 -14
rect 327 -15 328 -14
rect 328 -15 329 -14
rect 329 -15 330 -14
rect 330 -15 331 -14
rect 331 -15 332 -14
rect 332 -15 333 -14
rect 333 -15 334 -14
rect 334 -15 335 -14
rect 335 -15 336 -14
rect 336 -15 337 -14
rect 337 -15 338 -14
rect 338 -15 339 -14
rect 339 -15 340 -14
rect 340 -15 341 -14
rect 341 -15 342 -14
rect 342 -15 343 -14
rect 343 -15 344 -14
rect 344 -15 345 -14
rect 345 -15 346 -14
rect 346 -15 347 -14
rect 347 -15 348 -14
rect 348 -15 349 -14
rect 349 -15 350 -14
rect 350 -15 351 -14
rect 351 -15 352 -14
rect 352 -15 353 -14
rect 353 -15 354 -14
rect 354 -15 355 -14
rect 355 -15 356 -14
rect 356 -15 357 -14
rect 357 -15 358 -14
rect 358 -15 359 -14
rect 359 -15 360 -14
rect 360 -15 361 -14
rect 361 -15 362 -14
rect 362 -15 363 -14
rect 363 -15 364 -14
rect 364 -15 365 -14
rect 365 -15 366 -14
rect 366 -15 367 -14
rect 367 -15 368 -14
rect 368 -15 369 -14
rect 369 -15 370 -14
rect 370 -15 371 -14
rect 371 -15 372 -14
rect 372 -15 373 -14
rect 373 -15 374 -14
rect 374 -15 375 -14
rect 375 -15 376 -14
rect 376 -15 377 -14
rect 377 -15 378 -14
rect 378 -15 379 -14
rect 379 -15 380 -14
rect 380 -15 381 -14
rect 381 -15 382 -14
rect 382 -15 383 -14
rect 383 -15 384 -14
rect 384 -15 385 -14
rect 385 -15 386 -14
rect 386 -15 387 -14
rect 387 -15 388 -14
rect 388 -15 389 -14
rect 389 -15 390 -14
rect 390 -15 391 -14
rect 391 -15 392 -14
rect 392 -15 393 -14
rect 393 -15 394 -14
rect 394 -15 395 -14
rect 395 -15 396 -14
rect 396 -15 397 -14
rect 397 -15 398 -14
rect 398 -15 399 -14
rect 399 -15 400 -14
rect 400 -15 401 -14
rect 401 -15 402 -14
rect 402 -15 403 -14
rect 403 -15 404 -14
rect 404 -15 405 -14
rect 405 -15 406 -14
rect 406 -15 407 -14
rect 407 -15 408 -14
rect 408 -15 409 -14
rect 409 -15 410 -14
rect 410 -15 411 -14
rect 411 -15 412 -14
rect 412 -15 413 -14
rect 413 -15 414 -14
rect 414 -15 415 -14
rect 415 -15 416 -14
rect 416 -15 417 -14
rect 417 -15 418 -14
rect 418 -15 419 -14
rect 419 -15 420 -14
rect 420 -15 421 -14
rect 421 -15 422 -14
rect 422 -15 423 -14
rect 423 -15 424 -14
rect 424 -15 425 -14
rect 425 -15 426 -14
rect 426 -15 427 -14
rect 427 -15 428 -14
rect 428 -15 429 -14
rect 429 -15 430 -14
rect 430 -15 431 -14
rect 431 -15 432 -14
rect 432 -15 433 -14
rect 433 -15 434 -14
rect 434 -15 435 -14
rect 435 -15 436 -14
rect 436 -15 437 -14
rect 437 -15 438 -14
rect 438 -15 439 -14
rect 439 -15 440 -14
rect 440 -15 441 -14
rect 441 -15 442 -14
rect 442 -15 443 -14
rect 443 -15 444 -14
rect 444 -15 445 -14
rect 445 -15 446 -14
rect 446 -15 447 -14
rect 447 -15 448 -14
rect 448 -15 449 -14
rect 449 -15 450 -14
rect 450 -15 451 -14
rect 451 -15 452 -14
rect 452 -15 453 -14
rect 453 -15 454 -14
rect 454 -15 455 -14
rect 455 -15 456 -14
rect 456 -15 457 -14
rect 457 -15 458 -14
rect 458 -15 459 -14
rect 459 -15 460 -14
rect 460 -15 461 -14
rect 461 -15 462 -14
rect 462 -15 463 -14
rect 463 -15 464 -14
rect 464 -15 465 -14
rect 465 -15 466 -14
rect 466 -15 467 -14
rect 467 -15 468 -14
rect 468 -15 469 -14
rect 469 -15 470 -14
rect 470 -15 471 -14
rect 471 -15 472 -14
rect 472 -15 473 -14
rect 473 -15 474 -14
rect 474 -15 475 -14
rect 475 -15 476 -14
rect 476 -15 477 -14
rect 477 -15 478 -14
rect 478 -15 479 -14
rect 479 -15 480 -14
rect 2 -16 3 -15
rect 3 -16 4 -15
rect 4 -16 5 -15
rect 5 -16 6 -15
rect 6 -16 7 -15
rect 7 -16 8 -15
rect 8 -16 9 -15
rect 9 -16 10 -15
rect 10 -16 11 -15
rect 11 -16 12 -15
rect 21 -16 22 -15
rect 22 -16 23 -15
rect 23 -16 24 -15
rect 24 -16 25 -15
rect 25 -16 26 -15
rect 26 -16 27 -15
rect 27 -16 28 -15
rect 28 -16 29 -15
rect 29 -16 30 -15
rect 30 -16 31 -15
rect 31 -16 32 -15
rect 32 -16 33 -15
rect 33 -16 34 -15
rect 34 -16 35 -15
rect 35 -16 36 -15
rect 36 -16 37 -15
rect 37 -16 38 -15
rect 38 -16 39 -15
rect 39 -16 40 -15
rect 40 -16 41 -15
rect 41 -16 42 -15
rect 42 -16 43 -15
rect 43 -16 44 -15
rect 53 -16 54 -15
rect 54 -16 55 -15
rect 55 -16 56 -15
rect 56 -16 57 -15
rect 57 -16 58 -15
rect 58 -16 59 -15
rect 59 -16 60 -15
rect 60 -16 61 -15
rect 61 -16 62 -15
rect 62 -16 63 -15
rect 63 -16 64 -15
rect 64 -16 65 -15
rect 65 -16 66 -15
rect 66 -16 67 -15
rect 67 -16 68 -15
rect 68 -16 69 -15
rect 69 -16 70 -15
rect 70 -16 71 -15
rect 71 -16 72 -15
rect 72 -16 73 -15
rect 73 -16 74 -15
rect 74 -16 75 -15
rect 75 -16 76 -15
rect 85 -16 86 -15
rect 86 -16 87 -15
rect 87 -16 88 -15
rect 88 -16 89 -15
rect 89 -16 90 -15
rect 90 -16 91 -15
rect 91 -16 92 -15
rect 92 -16 93 -15
rect 93 -16 94 -15
rect 94 -16 95 -15
rect 95 -16 96 -15
rect 96 -16 97 -15
rect 97 -16 98 -15
rect 98 -16 99 -15
rect 99 -16 100 -15
rect 100 -16 101 -15
rect 101 -16 102 -15
rect 102 -16 103 -15
rect 103 -16 104 -15
rect 104 -16 105 -15
rect 105 -16 106 -15
rect 106 -16 107 -15
rect 107 -16 108 -15
rect 117 -16 118 -15
rect 118 -16 119 -15
rect 119 -16 120 -15
rect 120 -16 121 -15
rect 121 -16 122 -15
rect 122 -16 123 -15
rect 123 -16 124 -15
rect 124 -16 125 -15
rect 125 -16 126 -15
rect 126 -16 127 -15
rect 127 -16 128 -15
rect 128 -16 129 -15
rect 129 -16 130 -15
rect 130 -16 131 -15
rect 131 -16 132 -15
rect 132 -16 133 -15
rect 133 -16 134 -15
rect 134 -16 135 -15
rect 135 -16 136 -15
rect 136 -16 137 -15
rect 137 -16 138 -15
rect 138 -16 139 -15
rect 139 -16 140 -15
rect 149 -16 150 -15
rect 150 -16 151 -15
rect 151 -16 152 -15
rect 152 -16 153 -15
rect 153 -16 154 -15
rect 154 -16 155 -15
rect 155 -16 156 -15
rect 156 -16 157 -15
rect 157 -16 158 -15
rect 158 -16 159 -15
rect 159 -16 160 -15
rect 160 -16 161 -15
rect 161 -16 162 -15
rect 162 -16 163 -15
rect 163 -16 164 -15
rect 164 -16 165 -15
rect 165 -16 166 -15
rect 166 -16 167 -15
rect 167 -16 168 -15
rect 168 -16 169 -15
rect 169 -16 170 -15
rect 170 -16 171 -15
rect 171 -16 172 -15
rect 181 -16 182 -15
rect 182 -16 183 -15
rect 183 -16 184 -15
rect 184 -16 185 -15
rect 185 -16 186 -15
rect 186 -16 187 -15
rect 187 -16 188 -15
rect 188 -16 189 -15
rect 189 -16 190 -15
rect 190 -16 191 -15
rect 191 -16 192 -15
rect 192 -16 193 -15
rect 193 -16 194 -15
rect 194 -16 195 -15
rect 195 -16 196 -15
rect 196 -16 197 -15
rect 197 -16 198 -15
rect 198 -16 199 -15
rect 199 -16 200 -15
rect 200 -16 201 -15
rect 201 -16 202 -15
rect 202 -16 203 -15
rect 203 -16 204 -15
rect 204 -16 205 -15
rect 205 -16 206 -15
rect 206 -16 207 -15
rect 207 -16 208 -15
rect 208 -16 209 -15
rect 209 -16 210 -15
rect 210 -16 211 -15
rect 211 -16 212 -15
rect 212 -16 213 -15
rect 213 -16 214 -15
rect 214 -16 215 -15
rect 215 -16 216 -15
rect 216 -16 217 -15
rect 217 -16 218 -15
rect 218 -16 219 -15
rect 219 -16 220 -15
rect 220 -16 221 -15
rect 221 -16 222 -15
rect 222 -16 223 -15
rect 223 -16 224 -15
rect 224 -16 225 -15
rect 225 -16 226 -15
rect 226 -16 227 -15
rect 227 -16 228 -15
rect 228 -16 229 -15
rect 229 -16 230 -15
rect 230 -16 231 -15
rect 231 -16 232 -15
rect 232 -16 233 -15
rect 233 -16 234 -15
rect 234 -16 235 -15
rect 235 -16 236 -15
rect 236 -16 237 -15
rect 237 -16 238 -15
rect 238 -16 239 -15
rect 239 -16 240 -15
rect 240 -16 241 -15
rect 241 -16 242 -15
rect 242 -16 243 -15
rect 243 -16 244 -15
rect 244 -16 245 -15
rect 245 -16 246 -15
rect 246 -16 247 -15
rect 247 -16 248 -15
rect 248 -16 249 -15
rect 249 -16 250 -15
rect 250 -16 251 -15
rect 251 -16 252 -15
rect 252 -16 253 -15
rect 253 -16 254 -15
rect 254 -16 255 -15
rect 255 -16 256 -15
rect 256 -16 257 -15
rect 257 -16 258 -15
rect 258 -16 259 -15
rect 259 -16 260 -15
rect 260 -16 261 -15
rect 261 -16 262 -15
rect 262 -16 263 -15
rect 263 -16 264 -15
rect 264 -16 265 -15
rect 265 -16 266 -15
rect 266 -16 267 -15
rect 267 -16 268 -15
rect 268 -16 269 -15
rect 269 -16 270 -15
rect 270 -16 271 -15
rect 271 -16 272 -15
rect 272 -16 273 -15
rect 273 -16 274 -15
rect 274 -16 275 -15
rect 275 -16 276 -15
rect 276 -16 277 -15
rect 277 -16 278 -15
rect 278 -16 279 -15
rect 279 -16 280 -15
rect 280 -16 281 -15
rect 281 -16 282 -15
rect 282 -16 283 -15
rect 283 -16 284 -15
rect 284 -16 285 -15
rect 285 -16 286 -15
rect 286 -16 287 -15
rect 287 -16 288 -15
rect 288 -16 289 -15
rect 289 -16 290 -15
rect 290 -16 291 -15
rect 291 -16 292 -15
rect 292 -16 293 -15
rect 293 -16 294 -15
rect 294 -16 295 -15
rect 295 -16 296 -15
rect 296 -16 297 -15
rect 297 -16 298 -15
rect 298 -16 299 -15
rect 299 -16 300 -15
rect 300 -16 301 -15
rect 301 -16 302 -15
rect 302 -16 303 -15
rect 303 -16 304 -15
rect 304 -16 305 -15
rect 305 -16 306 -15
rect 306 -16 307 -15
rect 307 -16 308 -15
rect 308 -16 309 -15
rect 309 -16 310 -15
rect 310 -16 311 -15
rect 311 -16 312 -15
rect 312 -16 313 -15
rect 313 -16 314 -15
rect 314 -16 315 -15
rect 315 -16 316 -15
rect 316 -16 317 -15
rect 317 -16 318 -15
rect 318 -16 319 -15
rect 319 -16 320 -15
rect 320 -16 321 -15
rect 321 -16 322 -15
rect 322 -16 323 -15
rect 323 -16 324 -15
rect 324 -16 325 -15
rect 325 -16 326 -15
rect 326 -16 327 -15
rect 327 -16 328 -15
rect 328 -16 329 -15
rect 329 -16 330 -15
rect 330 -16 331 -15
rect 331 -16 332 -15
rect 332 -16 333 -15
rect 333 -16 334 -15
rect 334 -16 335 -15
rect 335 -16 336 -15
rect 336 -16 337 -15
rect 337 -16 338 -15
rect 338 -16 339 -15
rect 339 -16 340 -15
rect 340 -16 341 -15
rect 341 -16 342 -15
rect 342 -16 343 -15
rect 343 -16 344 -15
rect 344 -16 345 -15
rect 345 -16 346 -15
rect 346 -16 347 -15
rect 347 -16 348 -15
rect 348 -16 349 -15
rect 349 -16 350 -15
rect 350 -16 351 -15
rect 351 -16 352 -15
rect 352 -16 353 -15
rect 353 -16 354 -15
rect 354 -16 355 -15
rect 355 -16 356 -15
rect 356 -16 357 -15
rect 357 -16 358 -15
rect 358 -16 359 -15
rect 359 -16 360 -15
rect 360 -16 361 -15
rect 361 -16 362 -15
rect 362 -16 363 -15
rect 363 -16 364 -15
rect 364 -16 365 -15
rect 365 -16 366 -15
rect 366 -16 367 -15
rect 367 -16 368 -15
rect 368 -16 369 -15
rect 369 -16 370 -15
rect 370 -16 371 -15
rect 371 -16 372 -15
rect 372 -16 373 -15
rect 373 -16 374 -15
rect 374 -16 375 -15
rect 375 -16 376 -15
rect 376 -16 377 -15
rect 377 -16 378 -15
rect 378 -16 379 -15
rect 379 -16 380 -15
rect 380 -16 381 -15
rect 381 -16 382 -15
rect 382 -16 383 -15
rect 383 -16 384 -15
rect 384 -16 385 -15
rect 385 -16 386 -15
rect 386 -16 387 -15
rect 387 -16 388 -15
rect 388 -16 389 -15
rect 389 -16 390 -15
rect 390 -16 391 -15
rect 391 -16 392 -15
rect 392 -16 393 -15
rect 393 -16 394 -15
rect 394 -16 395 -15
rect 395 -16 396 -15
rect 396 -16 397 -15
rect 397 -16 398 -15
rect 398 -16 399 -15
rect 399 -16 400 -15
rect 400 -16 401 -15
rect 401 -16 402 -15
rect 402 -16 403 -15
rect 403 -16 404 -15
rect 404 -16 405 -15
rect 405 -16 406 -15
rect 406 -16 407 -15
rect 407 -16 408 -15
rect 408 -16 409 -15
rect 409 -16 410 -15
rect 410 -16 411 -15
rect 411 -16 412 -15
rect 412 -16 413 -15
rect 413 -16 414 -15
rect 414 -16 415 -15
rect 415 -16 416 -15
rect 416 -16 417 -15
rect 417 -16 418 -15
rect 418 -16 419 -15
rect 419 -16 420 -15
rect 420 -16 421 -15
rect 421 -16 422 -15
rect 422 -16 423 -15
rect 423 -16 424 -15
rect 424 -16 425 -15
rect 425 -16 426 -15
rect 426 -16 427 -15
rect 427 -16 428 -15
rect 428 -16 429 -15
rect 429 -16 430 -15
rect 430 -16 431 -15
rect 431 -16 432 -15
rect 432 -16 433 -15
rect 433 -16 434 -15
rect 434 -16 435 -15
rect 435 -16 436 -15
rect 436 -16 437 -15
rect 437 -16 438 -15
rect 438 -16 439 -15
rect 439 -16 440 -15
rect 440 -16 441 -15
rect 441 -16 442 -15
rect 442 -16 443 -15
rect 443 -16 444 -15
rect 444 -16 445 -15
rect 445 -16 446 -15
rect 446 -16 447 -15
rect 447 -16 448 -15
rect 448 -16 449 -15
rect 449 -16 450 -15
rect 450 -16 451 -15
rect 451 -16 452 -15
rect 452 -16 453 -15
rect 453 -16 454 -15
rect 454 -16 455 -15
rect 455 -16 456 -15
rect 456 -16 457 -15
rect 457 -16 458 -15
rect 458 -16 459 -15
rect 459 -16 460 -15
rect 460 -16 461 -15
rect 461 -16 462 -15
rect 462 -16 463 -15
rect 463 -16 464 -15
rect 464 -16 465 -15
rect 465 -16 466 -15
rect 466 -16 467 -15
rect 467 -16 468 -15
rect 468 -16 469 -15
rect 469 -16 470 -15
rect 470 -16 471 -15
rect 471 -16 472 -15
rect 472 -16 473 -15
rect 473 -16 474 -15
rect 474 -16 475 -15
rect 475 -16 476 -15
rect 476 -16 477 -15
rect 477 -16 478 -15
rect 478 -16 479 -15
rect 479 -16 480 -15
rect 2 -17 3 -16
rect 3 -17 4 -16
rect 4 -17 5 -16
rect 5 -17 6 -16
rect 6 -17 7 -16
rect 7 -17 8 -16
rect 8 -17 9 -16
rect 9 -17 10 -16
rect 10 -17 11 -16
rect 11 -17 12 -16
rect 21 -17 22 -16
rect 22 -17 23 -16
rect 23 -17 24 -16
rect 24 -17 25 -16
rect 25 -17 26 -16
rect 26 -17 27 -16
rect 27 -17 28 -16
rect 28 -17 29 -16
rect 29 -17 30 -16
rect 30 -17 31 -16
rect 31 -17 32 -16
rect 32 -17 33 -16
rect 33 -17 34 -16
rect 34 -17 35 -16
rect 35 -17 36 -16
rect 36 -17 37 -16
rect 37 -17 38 -16
rect 38 -17 39 -16
rect 39 -17 40 -16
rect 40 -17 41 -16
rect 41 -17 42 -16
rect 42 -17 43 -16
rect 43 -17 44 -16
rect 53 -17 54 -16
rect 54 -17 55 -16
rect 55 -17 56 -16
rect 56 -17 57 -16
rect 57 -17 58 -16
rect 58 -17 59 -16
rect 59 -17 60 -16
rect 60 -17 61 -16
rect 61 -17 62 -16
rect 62 -17 63 -16
rect 63 -17 64 -16
rect 64 -17 65 -16
rect 65 -17 66 -16
rect 66 -17 67 -16
rect 67 -17 68 -16
rect 68 -17 69 -16
rect 69 -17 70 -16
rect 70 -17 71 -16
rect 71 -17 72 -16
rect 72 -17 73 -16
rect 73 -17 74 -16
rect 74 -17 75 -16
rect 75 -17 76 -16
rect 85 -17 86 -16
rect 86 -17 87 -16
rect 87 -17 88 -16
rect 88 -17 89 -16
rect 89 -17 90 -16
rect 90 -17 91 -16
rect 91 -17 92 -16
rect 92 -17 93 -16
rect 93 -17 94 -16
rect 94 -17 95 -16
rect 95 -17 96 -16
rect 96 -17 97 -16
rect 97 -17 98 -16
rect 98 -17 99 -16
rect 99 -17 100 -16
rect 100 -17 101 -16
rect 101 -17 102 -16
rect 102 -17 103 -16
rect 103 -17 104 -16
rect 104 -17 105 -16
rect 105 -17 106 -16
rect 106 -17 107 -16
rect 107 -17 108 -16
rect 117 -17 118 -16
rect 118 -17 119 -16
rect 119 -17 120 -16
rect 120 -17 121 -16
rect 121 -17 122 -16
rect 122 -17 123 -16
rect 123 -17 124 -16
rect 124 -17 125 -16
rect 125 -17 126 -16
rect 126 -17 127 -16
rect 127 -17 128 -16
rect 128 -17 129 -16
rect 129 -17 130 -16
rect 130 -17 131 -16
rect 131 -17 132 -16
rect 132 -17 133 -16
rect 133 -17 134 -16
rect 134 -17 135 -16
rect 135 -17 136 -16
rect 136 -17 137 -16
rect 137 -17 138 -16
rect 138 -17 139 -16
rect 139 -17 140 -16
rect 149 -17 150 -16
rect 150 -17 151 -16
rect 151 -17 152 -16
rect 152 -17 153 -16
rect 153 -17 154 -16
rect 154 -17 155 -16
rect 155 -17 156 -16
rect 156 -17 157 -16
rect 157 -17 158 -16
rect 158 -17 159 -16
rect 159 -17 160 -16
rect 160 -17 161 -16
rect 161 -17 162 -16
rect 162 -17 163 -16
rect 163 -17 164 -16
rect 164 -17 165 -16
rect 165 -17 166 -16
rect 166 -17 167 -16
rect 167 -17 168 -16
rect 168 -17 169 -16
rect 169 -17 170 -16
rect 170 -17 171 -16
rect 171 -17 172 -16
rect 181 -17 182 -16
rect 182 -17 183 -16
rect 183 -17 184 -16
rect 184 -17 185 -16
rect 185 -17 186 -16
rect 186 -17 187 -16
rect 187 -17 188 -16
rect 188 -17 189 -16
rect 189 -17 190 -16
rect 190 -17 191 -16
rect 191 -17 192 -16
rect 192 -17 193 -16
rect 193 -17 194 -16
rect 194 -17 195 -16
rect 195 -17 196 -16
rect 196 -17 197 -16
rect 197 -17 198 -16
rect 198 -17 199 -16
rect 199 -17 200 -16
rect 200 -17 201 -16
rect 201 -17 202 -16
rect 202 -17 203 -16
rect 203 -17 204 -16
rect 204 -17 205 -16
rect 205 -17 206 -16
rect 206 -17 207 -16
rect 207 -17 208 -16
rect 208 -17 209 -16
rect 209 -17 210 -16
rect 210 -17 211 -16
rect 211 -17 212 -16
rect 212 -17 213 -16
rect 213 -17 214 -16
rect 214 -17 215 -16
rect 215 -17 216 -16
rect 216 -17 217 -16
rect 217 -17 218 -16
rect 218 -17 219 -16
rect 219 -17 220 -16
rect 220 -17 221 -16
rect 221 -17 222 -16
rect 222 -17 223 -16
rect 223 -17 224 -16
rect 224 -17 225 -16
rect 225 -17 226 -16
rect 226 -17 227 -16
rect 227 -17 228 -16
rect 228 -17 229 -16
rect 229 -17 230 -16
rect 230 -17 231 -16
rect 231 -17 232 -16
rect 232 -17 233 -16
rect 233 -17 234 -16
rect 234 -17 235 -16
rect 235 -17 236 -16
rect 236 -17 237 -16
rect 237 -17 238 -16
rect 238 -17 239 -16
rect 239 -17 240 -16
rect 240 -17 241 -16
rect 241 -17 242 -16
rect 242 -17 243 -16
rect 243 -17 244 -16
rect 244 -17 245 -16
rect 245 -17 246 -16
rect 246 -17 247 -16
rect 247 -17 248 -16
rect 248 -17 249 -16
rect 249 -17 250 -16
rect 250 -17 251 -16
rect 251 -17 252 -16
rect 252 -17 253 -16
rect 253 -17 254 -16
rect 254 -17 255 -16
rect 255 -17 256 -16
rect 256 -17 257 -16
rect 257 -17 258 -16
rect 258 -17 259 -16
rect 259 -17 260 -16
rect 260 -17 261 -16
rect 261 -17 262 -16
rect 262 -17 263 -16
rect 263 -17 264 -16
rect 264 -17 265 -16
rect 265 -17 266 -16
rect 266 -17 267 -16
rect 267 -17 268 -16
rect 268 -17 269 -16
rect 269 -17 270 -16
rect 270 -17 271 -16
rect 271 -17 272 -16
rect 272 -17 273 -16
rect 273 -17 274 -16
rect 274 -17 275 -16
rect 275 -17 276 -16
rect 276 -17 277 -16
rect 277 -17 278 -16
rect 278 -17 279 -16
rect 279 -17 280 -16
rect 280 -17 281 -16
rect 281 -17 282 -16
rect 282 -17 283 -16
rect 283 -17 284 -16
rect 284 -17 285 -16
rect 285 -17 286 -16
rect 286 -17 287 -16
rect 287 -17 288 -16
rect 288 -17 289 -16
rect 289 -17 290 -16
rect 290 -17 291 -16
rect 291 -17 292 -16
rect 292 -17 293 -16
rect 293 -17 294 -16
rect 294 -17 295 -16
rect 295 -17 296 -16
rect 296 -17 297 -16
rect 297 -17 298 -16
rect 298 -17 299 -16
rect 299 -17 300 -16
rect 300 -17 301 -16
rect 301 -17 302 -16
rect 302 -17 303 -16
rect 303 -17 304 -16
rect 304 -17 305 -16
rect 305 -17 306 -16
rect 306 -17 307 -16
rect 307 -17 308 -16
rect 308 -17 309 -16
rect 309 -17 310 -16
rect 310 -17 311 -16
rect 311 -17 312 -16
rect 312 -17 313 -16
rect 313 -17 314 -16
rect 314 -17 315 -16
rect 315 -17 316 -16
rect 316 -17 317 -16
rect 317 -17 318 -16
rect 318 -17 319 -16
rect 319 -17 320 -16
rect 320 -17 321 -16
rect 321 -17 322 -16
rect 322 -17 323 -16
rect 323 -17 324 -16
rect 324 -17 325 -16
rect 325 -17 326 -16
rect 326 -17 327 -16
rect 327 -17 328 -16
rect 328 -17 329 -16
rect 329 -17 330 -16
rect 330 -17 331 -16
rect 331 -17 332 -16
rect 332 -17 333 -16
rect 333 -17 334 -16
rect 334 -17 335 -16
rect 335 -17 336 -16
rect 336 -17 337 -16
rect 337 -17 338 -16
rect 338 -17 339 -16
rect 339 -17 340 -16
rect 340 -17 341 -16
rect 341 -17 342 -16
rect 342 -17 343 -16
rect 343 -17 344 -16
rect 344 -17 345 -16
rect 345 -17 346 -16
rect 346 -17 347 -16
rect 347 -17 348 -16
rect 348 -17 349 -16
rect 349 -17 350 -16
rect 350 -17 351 -16
rect 351 -17 352 -16
rect 352 -17 353 -16
rect 353 -17 354 -16
rect 354 -17 355 -16
rect 355 -17 356 -16
rect 356 -17 357 -16
rect 357 -17 358 -16
rect 358 -17 359 -16
rect 359 -17 360 -16
rect 360 -17 361 -16
rect 361 -17 362 -16
rect 362 -17 363 -16
rect 363 -17 364 -16
rect 364 -17 365 -16
rect 365 -17 366 -16
rect 366 -17 367 -16
rect 367 -17 368 -16
rect 368 -17 369 -16
rect 369 -17 370 -16
rect 370 -17 371 -16
rect 371 -17 372 -16
rect 372 -17 373 -16
rect 373 -17 374 -16
rect 374 -17 375 -16
rect 375 -17 376 -16
rect 376 -17 377 -16
rect 377 -17 378 -16
rect 378 -17 379 -16
rect 379 -17 380 -16
rect 380 -17 381 -16
rect 381 -17 382 -16
rect 382 -17 383 -16
rect 383 -17 384 -16
rect 384 -17 385 -16
rect 385 -17 386 -16
rect 386 -17 387 -16
rect 387 -17 388 -16
rect 388 -17 389 -16
rect 389 -17 390 -16
rect 390 -17 391 -16
rect 391 -17 392 -16
rect 392 -17 393 -16
rect 393 -17 394 -16
rect 394 -17 395 -16
rect 395 -17 396 -16
rect 396 -17 397 -16
rect 397 -17 398 -16
rect 398 -17 399 -16
rect 399 -17 400 -16
rect 400 -17 401 -16
rect 401 -17 402 -16
rect 402 -17 403 -16
rect 403 -17 404 -16
rect 404 -17 405 -16
rect 405 -17 406 -16
rect 406 -17 407 -16
rect 407 -17 408 -16
rect 408 -17 409 -16
rect 409 -17 410 -16
rect 410 -17 411 -16
rect 411 -17 412 -16
rect 412 -17 413 -16
rect 413 -17 414 -16
rect 414 -17 415 -16
rect 415 -17 416 -16
rect 416 -17 417 -16
rect 417 -17 418 -16
rect 418 -17 419 -16
rect 419 -17 420 -16
rect 420 -17 421 -16
rect 421 -17 422 -16
rect 422 -17 423 -16
rect 423 -17 424 -16
rect 424 -17 425 -16
rect 425 -17 426 -16
rect 426 -17 427 -16
rect 427 -17 428 -16
rect 428 -17 429 -16
rect 429 -17 430 -16
rect 430 -17 431 -16
rect 431 -17 432 -16
rect 432 -17 433 -16
rect 433 -17 434 -16
rect 434 -17 435 -16
rect 435 -17 436 -16
rect 436 -17 437 -16
rect 437 -17 438 -16
rect 438 -17 439 -16
rect 439 -17 440 -16
rect 440 -17 441 -16
rect 441 -17 442 -16
rect 442 -17 443 -16
rect 443 -17 444 -16
rect 444 -17 445 -16
rect 445 -17 446 -16
rect 446 -17 447 -16
rect 447 -17 448 -16
rect 448 -17 449 -16
rect 449 -17 450 -16
rect 450 -17 451 -16
rect 451 -17 452 -16
rect 452 -17 453 -16
rect 453 -17 454 -16
rect 454 -17 455 -16
rect 455 -17 456 -16
rect 456 -17 457 -16
rect 457 -17 458 -16
rect 458 -17 459 -16
rect 459 -17 460 -16
rect 460 -17 461 -16
rect 461 -17 462 -16
rect 462 -17 463 -16
rect 463 -17 464 -16
rect 464 -17 465 -16
rect 465 -17 466 -16
rect 466 -17 467 -16
rect 467 -17 468 -16
rect 468 -17 469 -16
rect 469 -17 470 -16
rect 470 -17 471 -16
rect 471 -17 472 -16
rect 472 -17 473 -16
rect 473 -17 474 -16
rect 474 -17 475 -16
rect 475 -17 476 -16
rect 476 -17 477 -16
rect 477 -17 478 -16
rect 478 -17 479 -16
rect 479 -17 480 -16
rect 2 -18 3 -17
rect 3 -18 4 -17
rect 4 -18 5 -17
rect 5 -18 6 -17
rect 6 -18 7 -17
rect 7 -18 8 -17
rect 8 -18 9 -17
rect 9 -18 10 -17
rect 10 -18 11 -17
rect 11 -18 12 -17
rect 16 -18 17 -17
rect 22 -18 23 -17
rect 23 -18 24 -17
rect 24 -18 25 -17
rect 25 -18 26 -17
rect 26 -18 27 -17
rect 27 -18 28 -17
rect 28 -18 29 -17
rect 29 -18 30 -17
rect 30 -18 31 -17
rect 31 -18 32 -17
rect 32 -18 33 -17
rect 33 -18 34 -17
rect 34 -18 35 -17
rect 35 -18 36 -17
rect 36 -18 37 -17
rect 37 -18 38 -17
rect 38 -18 39 -17
rect 39 -18 40 -17
rect 40 -18 41 -17
rect 41 -18 42 -17
rect 42 -18 43 -17
rect 43 -18 44 -17
rect 48 -18 49 -17
rect 54 -18 55 -17
rect 55 -18 56 -17
rect 56 -18 57 -17
rect 57 -18 58 -17
rect 58 -18 59 -17
rect 59 -18 60 -17
rect 60 -18 61 -17
rect 61 -18 62 -17
rect 62 -18 63 -17
rect 63 -18 64 -17
rect 64 -18 65 -17
rect 65 -18 66 -17
rect 66 -18 67 -17
rect 67 -18 68 -17
rect 68 -18 69 -17
rect 69 -18 70 -17
rect 70 -18 71 -17
rect 71 -18 72 -17
rect 72 -18 73 -17
rect 73 -18 74 -17
rect 74 -18 75 -17
rect 75 -18 76 -17
rect 80 -18 81 -17
rect 86 -18 87 -17
rect 87 -18 88 -17
rect 88 -18 89 -17
rect 89 -18 90 -17
rect 90 -18 91 -17
rect 91 -18 92 -17
rect 92 -18 93 -17
rect 93 -18 94 -17
rect 94 -18 95 -17
rect 95 -18 96 -17
rect 96 -18 97 -17
rect 97 -18 98 -17
rect 98 -18 99 -17
rect 99 -18 100 -17
rect 100 -18 101 -17
rect 101 -18 102 -17
rect 102 -18 103 -17
rect 103 -18 104 -17
rect 104 -18 105 -17
rect 105 -18 106 -17
rect 106 -18 107 -17
rect 107 -18 108 -17
rect 112 -18 113 -17
rect 118 -18 119 -17
rect 119 -18 120 -17
rect 120 -18 121 -17
rect 121 -18 122 -17
rect 122 -18 123 -17
rect 123 -18 124 -17
rect 124 -18 125 -17
rect 125 -18 126 -17
rect 126 -18 127 -17
rect 127 -18 128 -17
rect 128 -18 129 -17
rect 129 -18 130 -17
rect 130 -18 131 -17
rect 131 -18 132 -17
rect 132 -18 133 -17
rect 133 -18 134 -17
rect 134 -18 135 -17
rect 135 -18 136 -17
rect 136 -18 137 -17
rect 137 -18 138 -17
rect 138 -18 139 -17
rect 139 -18 140 -17
rect 144 -18 145 -17
rect 150 -18 151 -17
rect 151 -18 152 -17
rect 152 -18 153 -17
rect 153 -18 154 -17
rect 154 -18 155 -17
rect 155 -18 156 -17
rect 156 -18 157 -17
rect 157 -18 158 -17
rect 158 -18 159 -17
rect 159 -18 160 -17
rect 160 -18 161 -17
rect 161 -18 162 -17
rect 162 -18 163 -17
rect 163 -18 164 -17
rect 164 -18 165 -17
rect 165 -18 166 -17
rect 166 -18 167 -17
rect 167 -18 168 -17
rect 168 -18 169 -17
rect 169 -18 170 -17
rect 170 -18 171 -17
rect 171 -18 172 -17
rect 176 -18 177 -17
rect 182 -18 183 -17
rect 183 -18 184 -17
rect 184 -18 185 -17
rect 185 -18 186 -17
rect 186 -18 187 -17
rect 187 -18 188 -17
rect 188 -18 189 -17
rect 189 -18 190 -17
rect 190 -18 191 -17
rect 191 -18 192 -17
rect 2 -19 3 -18
rect 3 -19 4 -18
rect 4 -19 5 -18
rect 5 -19 6 -18
rect 6 -19 7 -18
rect 7 -19 8 -18
rect 8 -19 9 -18
rect 9 -19 10 -18
rect 10 -19 11 -18
rect 11 -19 12 -18
rect 14 -19 15 -18
rect 15 -19 16 -18
rect 16 -19 17 -18
rect 17 -19 18 -18
rect 18 -19 19 -18
rect 22 -19 23 -18
rect 23 -19 24 -18
rect 24 -19 25 -18
rect 25 -19 26 -18
rect 26 -19 27 -18
rect 27 -19 28 -18
rect 28 -19 29 -18
rect 29 -19 30 -18
rect 30 -19 31 -18
rect 31 -19 32 -18
rect 34 -19 35 -18
rect 35 -19 36 -18
rect 36 -19 37 -18
rect 37 -19 38 -18
rect 38 -19 39 -18
rect 39 -19 40 -18
rect 40 -19 41 -18
rect 41 -19 42 -18
rect 42 -19 43 -18
rect 43 -19 44 -18
rect 46 -19 47 -18
rect 47 -19 48 -18
rect 48 -19 49 -18
rect 49 -19 50 -18
rect 50 -19 51 -18
rect 54 -19 55 -18
rect 55 -19 56 -18
rect 56 -19 57 -18
rect 57 -19 58 -18
rect 58 -19 59 -18
rect 59 -19 60 -18
rect 60 -19 61 -18
rect 61 -19 62 -18
rect 62 -19 63 -18
rect 63 -19 64 -18
rect 66 -19 67 -18
rect 67 -19 68 -18
rect 68 -19 69 -18
rect 69 -19 70 -18
rect 70 -19 71 -18
rect 71 -19 72 -18
rect 72 -19 73 -18
rect 73 -19 74 -18
rect 74 -19 75 -18
rect 75 -19 76 -18
rect 78 -19 79 -18
rect 79 -19 80 -18
rect 80 -19 81 -18
rect 81 -19 82 -18
rect 82 -19 83 -18
rect 86 -19 87 -18
rect 87 -19 88 -18
rect 88 -19 89 -18
rect 89 -19 90 -18
rect 90 -19 91 -18
rect 91 -19 92 -18
rect 92 -19 93 -18
rect 93 -19 94 -18
rect 94 -19 95 -18
rect 95 -19 96 -18
rect 98 -19 99 -18
rect 99 -19 100 -18
rect 100 -19 101 -18
rect 101 -19 102 -18
rect 102 -19 103 -18
rect 103 -19 104 -18
rect 104 -19 105 -18
rect 105 -19 106 -18
rect 106 -19 107 -18
rect 107 -19 108 -18
rect 110 -19 111 -18
rect 111 -19 112 -18
rect 112 -19 113 -18
rect 113 -19 114 -18
rect 114 -19 115 -18
rect 118 -19 119 -18
rect 119 -19 120 -18
rect 120 -19 121 -18
rect 121 -19 122 -18
rect 122 -19 123 -18
rect 123 -19 124 -18
rect 124 -19 125 -18
rect 125 -19 126 -18
rect 126 -19 127 -18
rect 127 -19 128 -18
rect 130 -19 131 -18
rect 131 -19 132 -18
rect 132 -19 133 -18
rect 133 -19 134 -18
rect 134 -19 135 -18
rect 135 -19 136 -18
rect 136 -19 137 -18
rect 137 -19 138 -18
rect 138 -19 139 -18
rect 139 -19 140 -18
rect 142 -19 143 -18
rect 143 -19 144 -18
rect 144 -19 145 -18
rect 145 -19 146 -18
rect 146 -19 147 -18
rect 150 -19 151 -18
rect 151 -19 152 -18
rect 152 -19 153 -18
rect 153 -19 154 -18
rect 154 -19 155 -18
rect 155 -19 156 -18
rect 156 -19 157 -18
rect 157 -19 158 -18
rect 158 -19 159 -18
rect 159 -19 160 -18
rect 162 -19 163 -18
rect 163 -19 164 -18
rect 164 -19 165 -18
rect 165 -19 166 -18
rect 166 -19 167 -18
rect 167 -19 168 -18
rect 168 -19 169 -18
rect 169 -19 170 -18
rect 170 -19 171 -18
rect 171 -19 172 -18
rect 174 -19 175 -18
rect 175 -19 176 -18
rect 176 -19 177 -18
rect 177 -19 178 -18
rect 178 -19 179 -18
rect 182 -19 183 -18
rect 183 -19 184 -18
rect 184 -19 185 -18
rect 185 -19 186 -18
rect 186 -19 187 -18
rect 187 -19 188 -18
rect 188 -19 189 -18
rect 189 -19 190 -18
rect 190 -19 191 -18
rect 191 -19 192 -18
rect 2 -20 3 -19
rect 3 -20 4 -19
rect 4 -20 5 -19
rect 5 -20 6 -19
rect 6 -20 7 -19
rect 7 -20 8 -19
rect 8 -20 9 -19
rect 9 -20 10 -19
rect 10 -20 11 -19
rect 11 -20 12 -19
rect 12 -20 13 -19
rect 13 -20 14 -19
rect 14 -20 15 -19
rect 15 -20 16 -19
rect 16 -20 17 -19
rect 17 -20 18 -19
rect 18 -20 19 -19
rect 19 -20 20 -19
rect 20 -20 21 -19
rect 21 -20 22 -19
rect 22 -20 23 -19
rect 23 -20 24 -19
rect 24 -20 25 -19
rect 25 -20 26 -19
rect 26 -20 27 -19
rect 27 -20 28 -19
rect 28 -20 29 -19
rect 29 -20 30 -19
rect 30 -20 31 -19
rect 34 -20 35 -19
rect 35 -20 36 -19
rect 36 -20 37 -19
rect 37 -20 38 -19
rect 38 -20 39 -19
rect 39 -20 40 -19
rect 40 -20 41 -19
rect 41 -20 42 -19
rect 42 -20 43 -19
rect 43 -20 44 -19
rect 44 -20 45 -19
rect 45 -20 46 -19
rect 46 -20 47 -19
rect 47 -20 48 -19
rect 48 -20 49 -19
rect 49 -20 50 -19
rect 50 -20 51 -19
rect 51 -20 52 -19
rect 52 -20 53 -19
rect 53 -20 54 -19
rect 54 -20 55 -19
rect 55 -20 56 -19
rect 56 -20 57 -19
rect 57 -20 58 -19
rect 58 -20 59 -19
rect 59 -20 60 -19
rect 60 -20 61 -19
rect 61 -20 62 -19
rect 62 -20 63 -19
rect 66 -20 67 -19
rect 67 -20 68 -19
rect 68 -20 69 -19
rect 69 -20 70 -19
rect 70 -20 71 -19
rect 71 -20 72 -19
rect 72 -20 73 -19
rect 73 -20 74 -19
rect 74 -20 75 -19
rect 75 -20 76 -19
rect 76 -20 77 -19
rect 77 -20 78 -19
rect 78 -20 79 -19
rect 79 -20 80 -19
rect 80 -20 81 -19
rect 81 -20 82 -19
rect 82 -20 83 -19
rect 83 -20 84 -19
rect 84 -20 85 -19
rect 85 -20 86 -19
rect 86 -20 87 -19
rect 87 -20 88 -19
rect 88 -20 89 -19
rect 89 -20 90 -19
rect 90 -20 91 -19
rect 91 -20 92 -19
rect 92 -20 93 -19
rect 93 -20 94 -19
rect 94 -20 95 -19
rect 98 -20 99 -19
rect 99 -20 100 -19
rect 100 -20 101 -19
rect 101 -20 102 -19
rect 102 -20 103 -19
rect 103 -20 104 -19
rect 104 -20 105 -19
rect 105 -20 106 -19
rect 106 -20 107 -19
rect 107 -20 108 -19
rect 108 -20 109 -19
rect 109 -20 110 -19
rect 110 -20 111 -19
rect 111 -20 112 -19
rect 112 -20 113 -19
rect 113 -20 114 -19
rect 114 -20 115 -19
rect 115 -20 116 -19
rect 116 -20 117 -19
rect 117 -20 118 -19
rect 118 -20 119 -19
rect 119 -20 120 -19
rect 120 -20 121 -19
rect 121 -20 122 -19
rect 122 -20 123 -19
rect 123 -20 124 -19
rect 124 -20 125 -19
rect 125 -20 126 -19
rect 126 -20 127 -19
rect 130 -20 131 -19
rect 131 -20 132 -19
rect 132 -20 133 -19
rect 133 -20 134 -19
rect 134 -20 135 -19
rect 135 -20 136 -19
rect 136 -20 137 -19
rect 137 -20 138 -19
rect 138 -20 139 -19
rect 139 -20 140 -19
rect 140 -20 141 -19
rect 141 -20 142 -19
rect 142 -20 143 -19
rect 143 -20 144 -19
rect 144 -20 145 -19
rect 145 -20 146 -19
rect 146 -20 147 -19
rect 147 -20 148 -19
rect 148 -20 149 -19
rect 149 -20 150 -19
rect 150 -20 151 -19
rect 151 -20 152 -19
rect 152 -20 153 -19
rect 153 -20 154 -19
rect 154 -20 155 -19
rect 155 -20 156 -19
rect 156 -20 157 -19
rect 157 -20 158 -19
rect 158 -20 159 -19
rect 162 -20 163 -19
rect 163 -20 164 -19
rect 164 -20 165 -19
rect 165 -20 166 -19
rect 166 -20 167 -19
rect 167 -20 168 -19
rect 168 -20 169 -19
rect 169 -20 170 -19
rect 170 -20 171 -19
rect 171 -20 172 -19
rect 172 -20 173 -19
rect 173 -20 174 -19
rect 174 -20 175 -19
rect 175 -20 176 -19
rect 176 -20 177 -19
rect 177 -20 178 -19
rect 178 -20 179 -19
rect 179 -20 180 -19
rect 180 -20 181 -19
rect 181 -20 182 -19
rect 182 -20 183 -19
rect 183 -20 184 -19
rect 184 -20 185 -19
rect 185 -20 186 -19
rect 186 -20 187 -19
rect 187 -20 188 -19
rect 188 -20 189 -19
rect 189 -20 190 -19
rect 190 -20 191 -19
rect 191 -20 192 -19
rect 2 -21 3 -20
rect 3 -21 4 -20
rect 4 -21 5 -20
rect 5 -21 6 -20
rect 6 -21 7 -20
rect 7 -21 8 -20
rect 8 -21 9 -20
rect 9 -21 10 -20
rect 10 -21 11 -20
rect 11 -21 12 -20
rect 12 -21 13 -20
rect 13 -21 14 -20
rect 14 -21 15 -20
rect 15 -21 16 -20
rect 16 -21 17 -20
rect 17 -21 18 -20
rect 18 -21 19 -20
rect 19 -21 20 -20
rect 20 -21 21 -20
rect 21 -21 22 -20
rect 22 -21 23 -20
rect 23 -21 24 -20
rect 24 -21 25 -20
rect 25 -21 26 -20
rect 26 -21 27 -20
rect 27 -21 28 -20
rect 28 -21 29 -20
rect 29 -21 30 -20
rect 30 -21 31 -20
rect 34 -21 35 -20
rect 35 -21 36 -20
rect 36 -21 37 -20
rect 37 -21 38 -20
rect 38 -21 39 -20
rect 39 -21 40 -20
rect 40 -21 41 -20
rect 41 -21 42 -20
rect 42 -21 43 -20
rect 43 -21 44 -20
rect 44 -21 45 -20
rect 45 -21 46 -20
rect 46 -21 47 -20
rect 47 -21 48 -20
rect 48 -21 49 -20
rect 49 -21 50 -20
rect 50 -21 51 -20
rect 51 -21 52 -20
rect 52 -21 53 -20
rect 53 -21 54 -20
rect 54 -21 55 -20
rect 55 -21 56 -20
rect 56 -21 57 -20
rect 57 -21 58 -20
rect 58 -21 59 -20
rect 59 -21 60 -20
rect 60 -21 61 -20
rect 61 -21 62 -20
rect 62 -21 63 -20
rect 66 -21 67 -20
rect 67 -21 68 -20
rect 68 -21 69 -20
rect 69 -21 70 -20
rect 70 -21 71 -20
rect 71 -21 72 -20
rect 72 -21 73 -20
rect 73 -21 74 -20
rect 74 -21 75 -20
rect 75 -21 76 -20
rect 76 -21 77 -20
rect 77 -21 78 -20
rect 78 -21 79 -20
rect 79 -21 80 -20
rect 80 -21 81 -20
rect 81 -21 82 -20
rect 82 -21 83 -20
rect 83 -21 84 -20
rect 84 -21 85 -20
rect 85 -21 86 -20
rect 86 -21 87 -20
rect 87 -21 88 -20
rect 88 -21 89 -20
rect 89 -21 90 -20
rect 90 -21 91 -20
rect 91 -21 92 -20
rect 92 -21 93 -20
rect 93 -21 94 -20
rect 94 -21 95 -20
rect 98 -21 99 -20
rect 99 -21 100 -20
rect 100 -21 101 -20
rect 101 -21 102 -20
rect 102 -21 103 -20
rect 103 -21 104 -20
rect 104 -21 105 -20
rect 105 -21 106 -20
rect 106 -21 107 -20
rect 107 -21 108 -20
rect 108 -21 109 -20
rect 109 -21 110 -20
rect 110 -21 111 -20
rect 111 -21 112 -20
rect 112 -21 113 -20
rect 113 -21 114 -20
rect 114 -21 115 -20
rect 115 -21 116 -20
rect 116 -21 117 -20
rect 117 -21 118 -20
rect 118 -21 119 -20
rect 119 -21 120 -20
rect 120 -21 121 -20
rect 121 -21 122 -20
rect 122 -21 123 -20
rect 123 -21 124 -20
rect 124 -21 125 -20
rect 125 -21 126 -20
rect 126 -21 127 -20
rect 130 -21 131 -20
rect 131 -21 132 -20
rect 132 -21 133 -20
rect 133 -21 134 -20
rect 134 -21 135 -20
rect 135 -21 136 -20
rect 136 -21 137 -20
rect 137 -21 138 -20
rect 138 -21 139 -20
rect 139 -21 140 -20
rect 140 -21 141 -20
rect 141 -21 142 -20
rect 142 -21 143 -20
rect 143 -21 144 -20
rect 144 -21 145 -20
rect 145 -21 146 -20
rect 146 -21 147 -20
rect 147 -21 148 -20
rect 148 -21 149 -20
rect 149 -21 150 -20
rect 150 -21 151 -20
rect 151 -21 152 -20
rect 152 -21 153 -20
rect 153 -21 154 -20
rect 154 -21 155 -20
rect 155 -21 156 -20
rect 156 -21 157 -20
rect 157 -21 158 -20
rect 158 -21 159 -20
rect 162 -21 163 -20
rect 163 -21 164 -20
rect 164 -21 165 -20
rect 165 -21 166 -20
rect 166 -21 167 -20
rect 167 -21 168 -20
rect 168 -21 169 -20
rect 169 -21 170 -20
rect 170 -21 171 -20
rect 171 -21 172 -20
rect 172 -21 173 -20
rect 173 -21 174 -20
rect 174 -21 175 -20
rect 175 -21 176 -20
rect 176 -21 177 -20
rect 177 -21 178 -20
rect 178 -21 179 -20
rect 179 -21 180 -20
rect 180 -21 181 -20
rect 181 -21 182 -20
rect 182 -21 183 -20
rect 183 -21 184 -20
rect 184 -21 185 -20
rect 185 -21 186 -20
rect 186 -21 187 -20
rect 187 -21 188 -20
rect 188 -21 189 -20
rect 189 -21 190 -20
rect 190 -21 191 -20
rect 191 -21 192 -20
rect 2 -22 3 -21
rect 3 -22 4 -21
rect 4 -22 5 -21
rect 5 -22 6 -21
rect 6 -22 7 -21
rect 7 -22 8 -21
rect 8 -22 9 -21
rect 9 -22 10 -21
rect 10 -22 11 -21
rect 11 -22 12 -21
rect 12 -22 13 -21
rect 13 -22 14 -21
rect 14 -22 15 -21
rect 15 -22 16 -21
rect 16 -22 17 -21
rect 17 -22 18 -21
rect 18 -22 19 -21
rect 19 -22 20 -21
rect 20 -22 21 -21
rect 21 -22 22 -21
rect 22 -22 23 -21
rect 23 -22 24 -21
rect 24 -22 25 -21
rect 25 -22 26 -21
rect 26 -22 27 -21
rect 27 -22 28 -21
rect 28 -22 29 -21
rect 29 -22 30 -21
rect 30 -22 31 -21
rect 35 -22 36 -21
rect 36 -22 37 -21
rect 37 -22 38 -21
rect 38 -22 39 -21
rect 39 -22 40 -21
rect 40 -22 41 -21
rect 41 -22 42 -21
rect 42 -22 43 -21
rect 43 -22 44 -21
rect 44 -22 45 -21
rect 45 -22 46 -21
rect 46 -22 47 -21
rect 47 -22 48 -21
rect 48 -22 49 -21
rect 49 -22 50 -21
rect 50 -22 51 -21
rect 51 -22 52 -21
rect 52 -22 53 -21
rect 53 -22 54 -21
rect 54 -22 55 -21
rect 55 -22 56 -21
rect 56 -22 57 -21
rect 57 -22 58 -21
rect 58 -22 59 -21
rect 59 -22 60 -21
rect 60 -22 61 -21
rect 61 -22 62 -21
rect 62 -22 63 -21
rect 67 -22 68 -21
rect 68 -22 69 -21
rect 69 -22 70 -21
rect 70 -22 71 -21
rect 71 -22 72 -21
rect 72 -22 73 -21
rect 73 -22 74 -21
rect 74 -22 75 -21
rect 75 -22 76 -21
rect 76 -22 77 -21
rect 77 -22 78 -21
rect 78 -22 79 -21
rect 79 -22 80 -21
rect 80 -22 81 -21
rect 81 -22 82 -21
rect 82 -22 83 -21
rect 83 -22 84 -21
rect 84 -22 85 -21
rect 85 -22 86 -21
rect 86 -22 87 -21
rect 87 -22 88 -21
rect 88 -22 89 -21
rect 89 -22 90 -21
rect 90 -22 91 -21
rect 91 -22 92 -21
rect 92 -22 93 -21
rect 93 -22 94 -21
rect 94 -22 95 -21
rect 99 -22 100 -21
rect 100 -22 101 -21
rect 101 -22 102 -21
rect 102 -22 103 -21
rect 103 -22 104 -21
rect 104 -22 105 -21
rect 105 -22 106 -21
rect 106 -22 107 -21
rect 107 -22 108 -21
rect 108 -22 109 -21
rect 109 -22 110 -21
rect 110 -22 111 -21
rect 111 -22 112 -21
rect 112 -22 113 -21
rect 113 -22 114 -21
rect 114 -22 115 -21
rect 115 -22 116 -21
rect 116 -22 117 -21
rect 117 -22 118 -21
rect 118 -22 119 -21
rect 119 -22 120 -21
rect 120 -22 121 -21
rect 121 -22 122 -21
rect 122 -22 123 -21
rect 123 -22 124 -21
rect 124 -22 125 -21
rect 125 -22 126 -21
rect 126 -22 127 -21
rect 131 -22 132 -21
rect 132 -22 133 -21
rect 133 -22 134 -21
rect 134 -22 135 -21
rect 135 -22 136 -21
rect 136 -22 137 -21
rect 137 -22 138 -21
rect 138 -22 139 -21
rect 139 -22 140 -21
rect 140 -22 141 -21
rect 141 -22 142 -21
rect 142 -22 143 -21
rect 143 -22 144 -21
rect 144 -22 145 -21
rect 145 -22 146 -21
rect 146 -22 147 -21
rect 147 -22 148 -21
rect 148 -22 149 -21
rect 149 -22 150 -21
rect 150 -22 151 -21
rect 151 -22 152 -21
rect 152 -22 153 -21
rect 153 -22 154 -21
rect 154 -22 155 -21
rect 155 -22 156 -21
rect 156 -22 157 -21
rect 157 -22 158 -21
rect 158 -22 159 -21
rect 163 -22 164 -21
rect 164 -22 165 -21
rect 165 -22 166 -21
rect 166 -22 167 -21
rect 167 -22 168 -21
rect 168 -22 169 -21
rect 169 -22 170 -21
rect 170 -22 171 -21
rect 171 -22 172 -21
rect 172 -22 173 -21
rect 173 -22 174 -21
rect 174 -22 175 -21
rect 175 -22 176 -21
rect 176 -22 177 -21
rect 177 -22 178 -21
rect 178 -22 179 -21
rect 179 -22 180 -21
rect 180 -22 181 -21
rect 181 -22 182 -21
rect 182 -22 183 -21
rect 183 -22 184 -21
rect 184 -22 185 -21
rect 185 -22 186 -21
rect 186 -22 187 -21
rect 187 -22 188 -21
rect 188 -22 189 -21
rect 189 -22 190 -21
rect 190 -22 191 -21
rect 191 -22 192 -21
rect 2 -23 3 -22
rect 3 -23 4 -22
rect 4 -23 5 -22
rect 5 -23 6 -22
rect 6 -23 7 -22
rect 7 -23 8 -22
rect 8 -23 9 -22
rect 9 -23 10 -22
rect 10 -23 11 -22
rect 11 -23 12 -22
rect 12 -23 13 -22
rect 13 -23 14 -22
rect 14 -23 15 -22
rect 15 -23 16 -22
rect 16 -23 17 -22
rect 17 -23 18 -22
rect 18 -23 19 -22
rect 19 -23 20 -22
rect 20 -23 21 -22
rect 21 -23 22 -22
rect 22 -23 23 -22
rect 23 -23 24 -22
rect 24 -23 25 -22
rect 25 -23 26 -22
rect 26 -23 27 -22
rect 27 -23 28 -22
rect 28 -23 29 -22
rect 29 -23 30 -22
rect 35 -23 36 -22
rect 36 -23 37 -22
rect 37 -23 38 -22
rect 38 -23 39 -22
rect 39 -23 40 -22
rect 40 -23 41 -22
rect 41 -23 42 -22
rect 42 -23 43 -22
rect 43 -23 44 -22
rect 44 -23 45 -22
rect 45 -23 46 -22
rect 46 -23 47 -22
rect 47 -23 48 -22
rect 48 -23 49 -22
rect 49 -23 50 -22
rect 50 -23 51 -22
rect 51 -23 52 -22
rect 52 -23 53 -22
rect 53 -23 54 -22
rect 54 -23 55 -22
rect 55 -23 56 -22
rect 56 -23 57 -22
rect 57 -23 58 -22
rect 58 -23 59 -22
rect 59 -23 60 -22
rect 60 -23 61 -22
rect 61 -23 62 -22
rect 67 -23 68 -22
rect 68 -23 69 -22
rect 69 -23 70 -22
rect 70 -23 71 -22
rect 71 -23 72 -22
rect 72 -23 73 -22
rect 73 -23 74 -22
rect 74 -23 75 -22
rect 75 -23 76 -22
rect 76 -23 77 -22
rect 77 -23 78 -22
rect 78 -23 79 -22
rect 79 -23 80 -22
rect 80 -23 81 -22
rect 81 -23 82 -22
rect 82 -23 83 -22
rect 83 -23 84 -22
rect 84 -23 85 -22
rect 85 -23 86 -22
rect 86 -23 87 -22
rect 87 -23 88 -22
rect 88 -23 89 -22
rect 89 -23 90 -22
rect 90 -23 91 -22
rect 91 -23 92 -22
rect 92 -23 93 -22
rect 93 -23 94 -22
rect 99 -23 100 -22
rect 100 -23 101 -22
rect 101 -23 102 -22
rect 102 -23 103 -22
rect 103 -23 104 -22
rect 104 -23 105 -22
rect 105 -23 106 -22
rect 106 -23 107 -22
rect 107 -23 108 -22
rect 108 -23 109 -22
rect 109 -23 110 -22
rect 110 -23 111 -22
rect 111 -23 112 -22
rect 112 -23 113 -22
rect 113 -23 114 -22
rect 114 -23 115 -22
rect 115 -23 116 -22
rect 116 -23 117 -22
rect 117 -23 118 -22
rect 118 -23 119 -22
rect 119 -23 120 -22
rect 120 -23 121 -22
rect 121 -23 122 -22
rect 122 -23 123 -22
rect 123 -23 124 -22
rect 124 -23 125 -22
rect 125 -23 126 -22
rect 131 -23 132 -22
rect 132 -23 133 -22
rect 133 -23 134 -22
rect 134 -23 135 -22
rect 135 -23 136 -22
rect 136 -23 137 -22
rect 137 -23 138 -22
rect 138 -23 139 -22
rect 139 -23 140 -22
rect 140 -23 141 -22
rect 141 -23 142 -22
rect 142 -23 143 -22
rect 143 -23 144 -22
rect 144 -23 145 -22
rect 145 -23 146 -22
rect 146 -23 147 -22
rect 147 -23 148 -22
rect 148 -23 149 -22
rect 149 -23 150 -22
rect 150 -23 151 -22
rect 151 -23 152 -22
rect 152 -23 153 -22
rect 153 -23 154 -22
rect 154 -23 155 -22
rect 155 -23 156 -22
rect 156 -23 157 -22
rect 157 -23 158 -22
rect 163 -23 164 -22
rect 164 -23 165 -22
rect 165 -23 166 -22
rect 166 -23 167 -22
rect 167 -23 168 -22
rect 168 -23 169 -22
rect 169 -23 170 -22
rect 170 -23 171 -22
rect 171 -23 172 -22
rect 172 -23 173 -22
rect 173 -23 174 -22
rect 174 -23 175 -22
rect 175 -23 176 -22
rect 176 -23 177 -22
rect 177 -23 178 -22
rect 178 -23 179 -22
rect 179 -23 180 -22
rect 180 -23 181 -22
rect 181 -23 182 -22
rect 182 -23 183 -22
rect 183 -23 184 -22
rect 184 -23 185 -22
rect 185 -23 186 -22
rect 186 -23 187 -22
rect 187 -23 188 -22
rect 188 -23 189 -22
rect 189 -23 190 -22
rect 190 -23 191 -22
rect 191 -23 192 -22
rect 2 -24 3 -23
rect 3 -24 4 -23
rect 4 -24 5 -23
rect 5 -24 6 -23
rect 6 -24 7 -23
rect 7 -24 8 -23
rect 8 -24 9 -23
rect 9 -24 10 -23
rect 10 -24 11 -23
rect 11 -24 12 -23
rect 12 -24 13 -23
rect 13 -24 14 -23
rect 14 -24 15 -23
rect 15 -24 16 -23
rect 16 -24 17 -23
rect 17 -24 18 -23
rect 18 -24 19 -23
rect 19 -24 20 -23
rect 20 -24 21 -23
rect 21 -24 22 -23
rect 22 -24 23 -23
rect 23 -24 24 -23
rect 24 -24 25 -23
rect 41 -24 42 -23
rect 42 -24 43 -23
rect 43 -24 44 -23
rect 44 -24 45 -23
rect 45 -24 46 -23
rect 46 -24 47 -23
rect 47 -24 48 -23
rect 48 -24 49 -23
rect 49 -24 50 -23
rect 50 -24 51 -23
rect 51 -24 52 -23
rect 52 -24 53 -23
rect 53 -24 54 -23
rect 54 -24 55 -23
rect 55 -24 56 -23
rect 56 -24 57 -23
rect 73 -24 74 -23
rect 74 -24 75 -23
rect 75 -24 76 -23
rect 76 -24 77 -23
rect 77 -24 78 -23
rect 78 -24 79 -23
rect 79 -24 80 -23
rect 80 -24 81 -23
rect 81 -24 82 -23
rect 82 -24 83 -23
rect 83 -24 84 -23
rect 84 -24 85 -23
rect 85 -24 86 -23
rect 86 -24 87 -23
rect 87 -24 88 -23
rect 88 -24 89 -23
rect 105 -24 106 -23
rect 106 -24 107 -23
rect 107 -24 108 -23
rect 108 -24 109 -23
rect 109 -24 110 -23
rect 110 -24 111 -23
rect 111 -24 112 -23
rect 112 -24 113 -23
rect 113 -24 114 -23
rect 114 -24 115 -23
rect 115 -24 116 -23
rect 116 -24 117 -23
rect 117 -24 118 -23
rect 118 -24 119 -23
rect 119 -24 120 -23
rect 120 -24 121 -23
rect 137 -24 138 -23
rect 138 -24 139 -23
rect 139 -24 140 -23
rect 140 -24 141 -23
rect 141 -24 142 -23
rect 142 -24 143 -23
rect 143 -24 144 -23
rect 144 -24 145 -23
rect 145 -24 146 -23
rect 146 -24 147 -23
rect 147 -24 148 -23
rect 148 -24 149 -23
rect 149 -24 150 -23
rect 150 -24 151 -23
rect 151 -24 152 -23
rect 152 -24 153 -23
rect 169 -24 170 -23
rect 170 -24 171 -23
rect 171 -24 172 -23
rect 172 -24 173 -23
rect 173 -24 174 -23
rect 174 -24 175 -23
rect 175 -24 176 -23
rect 176 -24 177 -23
rect 177 -24 178 -23
rect 178 -24 179 -23
rect 179 -24 180 -23
rect 180 -24 181 -23
rect 181 -24 182 -23
rect 182 -24 183 -23
rect 183 -24 184 -23
rect 184 -24 185 -23
rect 185 -24 186 -23
rect 186 -24 187 -23
rect 187 -24 188 -23
rect 188 -24 189 -23
rect 189 -24 190 -23
rect 190 -24 191 -23
rect 191 -24 192 -23
rect 2 -25 3 -24
rect 3 -25 4 -24
rect 4 -25 5 -24
rect 5 -25 6 -24
rect 6 -25 7 -24
rect 7 -25 8 -24
rect 8 -25 9 -24
rect 9 -25 10 -24
rect 10 -25 11 -24
rect 11 -25 12 -24
rect 12 -25 13 -24
rect 13 -25 14 -24
rect 14 -25 15 -24
rect 15 -25 16 -24
rect 16 -25 17 -24
rect 17 -25 18 -24
rect 18 -25 19 -24
rect 19 -25 20 -24
rect 20 -25 21 -24
rect 21 -25 22 -24
rect 22 -25 23 -24
rect 23 -25 24 -24
rect 24 -25 25 -24
rect 41 -25 42 -24
rect 42 -25 43 -24
rect 43 -25 44 -24
rect 44 -25 45 -24
rect 45 -25 46 -24
rect 46 -25 47 -24
rect 47 -25 48 -24
rect 48 -25 49 -24
rect 49 -25 50 -24
rect 50 -25 51 -24
rect 51 -25 52 -24
rect 52 -25 53 -24
rect 53 -25 54 -24
rect 54 -25 55 -24
rect 55 -25 56 -24
rect 56 -25 57 -24
rect 73 -25 74 -24
rect 74 -25 75 -24
rect 75 -25 76 -24
rect 76 -25 77 -24
rect 77 -25 78 -24
rect 78 -25 79 -24
rect 79 -25 80 -24
rect 80 -25 81 -24
rect 81 -25 82 -24
rect 82 -25 83 -24
rect 83 -25 84 -24
rect 84 -25 85 -24
rect 85 -25 86 -24
rect 86 -25 87 -24
rect 87 -25 88 -24
rect 88 -25 89 -24
rect 105 -25 106 -24
rect 106 -25 107 -24
rect 107 -25 108 -24
rect 108 -25 109 -24
rect 109 -25 110 -24
rect 110 -25 111 -24
rect 111 -25 112 -24
rect 112 -25 113 -24
rect 113 -25 114 -24
rect 114 -25 115 -24
rect 115 -25 116 -24
rect 116 -25 117 -24
rect 117 -25 118 -24
rect 118 -25 119 -24
rect 119 -25 120 -24
rect 120 -25 121 -24
rect 137 -25 138 -24
rect 138 -25 139 -24
rect 139 -25 140 -24
rect 140 -25 141 -24
rect 141 -25 142 -24
rect 142 -25 143 -24
rect 143 -25 144 -24
rect 144 -25 145 -24
rect 145 -25 146 -24
rect 146 -25 147 -24
rect 147 -25 148 -24
rect 148 -25 149 -24
rect 149 -25 150 -24
rect 150 -25 151 -24
rect 151 -25 152 -24
rect 152 -25 153 -24
rect 169 -25 170 -24
rect 170 -25 171 -24
rect 171 -25 172 -24
rect 172 -25 173 -24
rect 173 -25 174 -24
rect 174 -25 175 -24
rect 175 -25 176 -24
rect 176 -25 177 -24
rect 177 -25 178 -24
rect 178 -25 179 -24
rect 179 -25 180 -24
rect 180 -25 181 -24
rect 181 -25 182 -24
rect 182 -25 183 -24
rect 183 -25 184 -24
rect 184 -25 185 -24
rect 185 -25 186 -24
rect 186 -25 187 -24
rect 187 -25 188 -24
rect 188 -25 189 -24
rect 189 -25 190 -24
rect 190 -25 191 -24
rect 191 -25 192 -24
rect 2 -26 3 -25
rect 3 -26 4 -25
rect 4 -26 5 -25
rect 5 -26 6 -25
rect 6 -26 7 -25
rect 7 -26 8 -25
rect 8 -26 9 -25
rect 9 -26 10 -25
rect 10 -26 11 -25
rect 11 -26 12 -25
rect 12 -26 13 -25
rect 13 -26 14 -25
rect 14 -26 15 -25
rect 15 -26 16 -25
rect 16 -26 17 -25
rect 17 -26 18 -25
rect 18 -26 19 -25
rect 19 -26 20 -25
rect 20 -26 21 -25
rect 21 -26 22 -25
rect 22 -26 23 -25
rect 23 -26 24 -25
rect 24 -26 25 -25
rect 25 -26 26 -25
rect 40 -26 41 -25
rect 41 -26 42 -25
rect 42 -26 43 -25
rect 43 -26 44 -25
rect 44 -26 45 -25
rect 45 -26 46 -25
rect 46 -26 47 -25
rect 47 -26 48 -25
rect 48 -26 49 -25
rect 49 -26 50 -25
rect 50 -26 51 -25
rect 51 -26 52 -25
rect 52 -26 53 -25
rect 53 -26 54 -25
rect 54 -26 55 -25
rect 55 -26 56 -25
rect 56 -26 57 -25
rect 57 -26 58 -25
rect 72 -26 73 -25
rect 73 -26 74 -25
rect 74 -26 75 -25
rect 75 -26 76 -25
rect 76 -26 77 -25
rect 77 -26 78 -25
rect 78 -26 79 -25
rect 79 -26 80 -25
rect 80 -26 81 -25
rect 81 -26 82 -25
rect 82 -26 83 -25
rect 83 -26 84 -25
rect 84 -26 85 -25
rect 85 -26 86 -25
rect 86 -26 87 -25
rect 87 -26 88 -25
rect 88 -26 89 -25
rect 89 -26 90 -25
rect 104 -26 105 -25
rect 105 -26 106 -25
rect 106 -26 107 -25
rect 107 -26 108 -25
rect 108 -26 109 -25
rect 109 -26 110 -25
rect 110 -26 111 -25
rect 111 -26 112 -25
rect 112 -26 113 -25
rect 113 -26 114 -25
rect 114 -26 115 -25
rect 115 -26 116 -25
rect 116 -26 117 -25
rect 117 -26 118 -25
rect 118 -26 119 -25
rect 119 -26 120 -25
rect 120 -26 121 -25
rect 121 -26 122 -25
rect 136 -26 137 -25
rect 137 -26 138 -25
rect 138 -26 139 -25
rect 139 -26 140 -25
rect 140 -26 141 -25
rect 141 -26 142 -25
rect 142 -26 143 -25
rect 143 -26 144 -25
rect 144 -26 145 -25
rect 145 -26 146 -25
rect 146 -26 147 -25
rect 147 -26 148 -25
rect 148 -26 149 -25
rect 149 -26 150 -25
rect 150 -26 151 -25
rect 151 -26 152 -25
rect 152 -26 153 -25
rect 153 -26 154 -25
rect 168 -26 169 -25
rect 169 -26 170 -25
rect 170 -26 171 -25
rect 171 -26 172 -25
rect 172 -26 173 -25
rect 173 -26 174 -25
rect 174 -26 175 -25
rect 175 -26 176 -25
rect 176 -26 177 -25
rect 177 -26 178 -25
rect 178 -26 179 -25
rect 179 -26 180 -25
rect 180 -26 181 -25
rect 181 -26 182 -25
rect 182 -26 183 -25
rect 183 -26 184 -25
rect 184 -26 185 -25
rect 185 -26 186 -25
rect 186 -26 187 -25
rect 187 -26 188 -25
rect 188 -26 189 -25
rect 189 -26 190 -25
rect 190 -26 191 -25
rect 191 -26 192 -25
rect 2 -27 3 -26
rect 3 -27 4 -26
rect 4 -27 5 -26
rect 5 -27 6 -26
rect 6 -27 7 -26
rect 7 -27 8 -26
rect 8 -27 9 -26
rect 9 -27 10 -26
rect 10 -27 11 -26
rect 11 -27 12 -26
rect 12 -27 13 -26
rect 13 -27 14 -26
rect 14 -27 15 -26
rect 15 -27 16 -26
rect 16 -27 17 -26
rect 17 -27 18 -26
rect 18 -27 19 -26
rect 19 -27 20 -26
rect 20 -27 21 -26
rect 21 -27 22 -26
rect 22 -27 23 -26
rect 23 -27 24 -26
rect 24 -27 25 -26
rect 25 -27 26 -26
rect 26 -27 27 -26
rect 38 -27 39 -26
rect 39 -27 40 -26
rect 40 -27 41 -26
rect 41 -27 42 -26
rect 42 -27 43 -26
rect 43 -27 44 -26
rect 44 -27 45 -26
rect 45 -27 46 -26
rect 46 -27 47 -26
rect 47 -27 48 -26
rect 48 -27 49 -26
rect 49 -27 50 -26
rect 50 -27 51 -26
rect 51 -27 52 -26
rect 52 -27 53 -26
rect 53 -27 54 -26
rect 54 -27 55 -26
rect 55 -27 56 -26
rect 56 -27 57 -26
rect 57 -27 58 -26
rect 58 -27 59 -26
rect 70 -27 71 -26
rect 71 -27 72 -26
rect 72 -27 73 -26
rect 73 -27 74 -26
rect 74 -27 75 -26
rect 75 -27 76 -26
rect 76 -27 77 -26
rect 77 -27 78 -26
rect 78 -27 79 -26
rect 79 -27 80 -26
rect 80 -27 81 -26
rect 81 -27 82 -26
rect 82 -27 83 -26
rect 83 -27 84 -26
rect 84 -27 85 -26
rect 85 -27 86 -26
rect 86 -27 87 -26
rect 87 -27 88 -26
rect 88 -27 89 -26
rect 89 -27 90 -26
rect 90 -27 91 -26
rect 102 -27 103 -26
rect 103 -27 104 -26
rect 104 -27 105 -26
rect 105 -27 106 -26
rect 106 -27 107 -26
rect 107 -27 108 -26
rect 108 -27 109 -26
rect 109 -27 110 -26
rect 110 -27 111 -26
rect 111 -27 112 -26
rect 112 -27 113 -26
rect 113 -27 114 -26
rect 114 -27 115 -26
rect 115 -27 116 -26
rect 116 -27 117 -26
rect 117 -27 118 -26
rect 118 -27 119 -26
rect 119 -27 120 -26
rect 120 -27 121 -26
rect 121 -27 122 -26
rect 122 -27 123 -26
rect 134 -27 135 -26
rect 135 -27 136 -26
rect 136 -27 137 -26
rect 137 -27 138 -26
rect 138 -27 139 -26
rect 139 -27 140 -26
rect 140 -27 141 -26
rect 141 -27 142 -26
rect 142 -27 143 -26
rect 143 -27 144 -26
rect 144 -27 145 -26
rect 145 -27 146 -26
rect 146 -27 147 -26
rect 147 -27 148 -26
rect 148 -27 149 -26
rect 149 -27 150 -26
rect 150 -27 151 -26
rect 151 -27 152 -26
rect 152 -27 153 -26
rect 153 -27 154 -26
rect 154 -27 155 -26
rect 166 -27 167 -26
rect 167 -27 168 -26
rect 168 -27 169 -26
rect 169 -27 170 -26
rect 170 -27 171 -26
rect 171 -27 172 -26
rect 172 -27 173 -26
rect 173 -27 174 -26
rect 174 -27 175 -26
rect 175 -27 176 -26
rect 176 -27 177 -26
rect 177 -27 178 -26
rect 178 -27 179 -26
rect 179 -27 180 -26
rect 180 -27 181 -26
rect 181 -27 182 -26
rect 182 -27 183 -26
rect 183 -27 184 -26
rect 184 -27 185 -26
rect 185 -27 186 -26
rect 186 -27 187 -26
rect 187 -27 188 -26
rect 188 -27 189 -26
rect 189 -27 190 -26
rect 190 -27 191 -26
rect 191 -27 192 -26
rect 2 -28 3 -27
rect 3 -28 4 -27
rect 4 -28 5 -27
rect 5 -28 6 -27
rect 6 -28 7 -27
rect 7 -28 8 -27
rect 8 -28 9 -27
rect 9 -28 10 -27
rect 10 -28 11 -27
rect 11 -28 12 -27
rect 12 -28 13 -27
rect 13 -28 14 -27
rect 14 -28 15 -27
rect 15 -28 16 -27
rect 16 -28 17 -27
rect 17 -28 18 -27
rect 18 -28 19 -27
rect 19 -28 20 -27
rect 20 -28 21 -27
rect 21 -28 22 -27
rect 22 -28 23 -27
rect 23 -28 24 -27
rect 24 -28 25 -27
rect 25 -28 26 -27
rect 26 -28 27 -27
rect 27 -28 28 -27
rect 37 -28 38 -27
rect 38 -28 39 -27
rect 39 -28 40 -27
rect 40 -28 41 -27
rect 41 -28 42 -27
rect 42 -28 43 -27
rect 43 -28 44 -27
rect 44 -28 45 -27
rect 45 -28 46 -27
rect 46 -28 47 -27
rect 47 -28 48 -27
rect 48 -28 49 -27
rect 49 -28 50 -27
rect 50 -28 51 -27
rect 51 -28 52 -27
rect 52 -28 53 -27
rect 53 -28 54 -27
rect 54 -28 55 -27
rect 55 -28 56 -27
rect 56 -28 57 -27
rect 57 -28 58 -27
rect 58 -28 59 -27
rect 59 -28 60 -27
rect 69 -28 70 -27
rect 70 -28 71 -27
rect 71 -28 72 -27
rect 72 -28 73 -27
rect 73 -28 74 -27
rect 74 -28 75 -27
rect 75 -28 76 -27
rect 76 -28 77 -27
rect 77 -28 78 -27
rect 78 -28 79 -27
rect 79 -28 80 -27
rect 80 -28 81 -27
rect 81 -28 82 -27
rect 82 -28 83 -27
rect 83 -28 84 -27
rect 84 -28 85 -27
rect 85 -28 86 -27
rect 86 -28 87 -27
rect 87 -28 88 -27
rect 88 -28 89 -27
rect 89 -28 90 -27
rect 90 -28 91 -27
rect 91 -28 92 -27
rect 101 -28 102 -27
rect 102 -28 103 -27
rect 103 -28 104 -27
rect 104 -28 105 -27
rect 105 -28 106 -27
rect 106 -28 107 -27
rect 107 -28 108 -27
rect 108 -28 109 -27
rect 109 -28 110 -27
rect 110 -28 111 -27
rect 111 -28 112 -27
rect 112 -28 113 -27
rect 113 -28 114 -27
rect 114 -28 115 -27
rect 115 -28 116 -27
rect 116 -28 117 -27
rect 117 -28 118 -27
rect 118 -28 119 -27
rect 119 -28 120 -27
rect 120 -28 121 -27
rect 121 -28 122 -27
rect 122 -28 123 -27
rect 123 -28 124 -27
rect 133 -28 134 -27
rect 134 -28 135 -27
rect 135 -28 136 -27
rect 136 -28 137 -27
rect 137 -28 138 -27
rect 138 -28 139 -27
rect 139 -28 140 -27
rect 140 -28 141 -27
rect 141 -28 142 -27
rect 142 -28 143 -27
rect 143 -28 144 -27
rect 144 -28 145 -27
rect 145 -28 146 -27
rect 146 -28 147 -27
rect 147 -28 148 -27
rect 148 -28 149 -27
rect 149 -28 150 -27
rect 150 -28 151 -27
rect 151 -28 152 -27
rect 152 -28 153 -27
rect 153 -28 154 -27
rect 154 -28 155 -27
rect 155 -28 156 -27
rect 165 -28 166 -27
rect 166 -28 167 -27
rect 167 -28 168 -27
rect 168 -28 169 -27
rect 169 -28 170 -27
rect 170 -28 171 -27
rect 171 -28 172 -27
rect 172 -28 173 -27
rect 173 -28 174 -27
rect 174 -28 175 -27
rect 175 -28 176 -27
rect 176 -28 177 -27
rect 177 -28 178 -27
rect 178 -28 179 -27
rect 179 -28 180 -27
rect 180 -28 181 -27
rect 181 -28 182 -27
rect 182 -28 183 -27
rect 183 -28 184 -27
rect 184 -28 185 -27
rect 185 -28 186 -27
rect 186 -28 187 -27
rect 187 -28 188 -27
rect 188 -28 189 -27
rect 189 -28 190 -27
rect 190 -28 191 -27
rect 191 -28 192 -27
rect 2 -29 3 -28
rect 3 -29 4 -28
rect 4 -29 5 -28
rect 5 -29 6 -28
rect 6 -29 7 -28
rect 7 -29 8 -28
rect 8 -29 9 -28
rect 9 -29 10 -28
rect 10 -29 11 -28
rect 11 -29 12 -28
rect 12 -29 13 -28
rect 13 -29 14 -28
rect 14 -29 15 -28
rect 15 -29 16 -28
rect 16 -29 17 -28
rect 17 -29 18 -28
rect 18 -29 19 -28
rect 19 -29 20 -28
rect 20 -29 21 -28
rect 21 -29 22 -28
rect 22 -29 23 -28
rect 23 -29 24 -28
rect 24 -29 25 -28
rect 25 -29 26 -28
rect 26 -29 27 -28
rect 27 -29 28 -28
rect 37 -29 38 -28
rect 38 -29 39 -28
rect 39 -29 40 -28
rect 40 -29 41 -28
rect 41 -29 42 -28
rect 42 -29 43 -28
rect 43 -29 44 -28
rect 44 -29 45 -28
rect 45 -29 46 -28
rect 46 -29 47 -28
rect 47 -29 48 -28
rect 48 -29 49 -28
rect 49 -29 50 -28
rect 50 -29 51 -28
rect 51 -29 52 -28
rect 52 -29 53 -28
rect 53 -29 54 -28
rect 54 -29 55 -28
rect 55 -29 56 -28
rect 56 -29 57 -28
rect 57 -29 58 -28
rect 58 -29 59 -28
rect 59 -29 60 -28
rect 69 -29 70 -28
rect 70 -29 71 -28
rect 71 -29 72 -28
rect 72 -29 73 -28
rect 73 -29 74 -28
rect 74 -29 75 -28
rect 75 -29 76 -28
rect 76 -29 77 -28
rect 77 -29 78 -28
rect 78 -29 79 -28
rect 79 -29 80 -28
rect 80 -29 81 -28
rect 81 -29 82 -28
rect 82 -29 83 -28
rect 83 -29 84 -28
rect 84 -29 85 -28
rect 85 -29 86 -28
rect 86 -29 87 -28
rect 87 -29 88 -28
rect 88 -29 89 -28
rect 89 -29 90 -28
rect 90 -29 91 -28
rect 91 -29 92 -28
rect 101 -29 102 -28
rect 102 -29 103 -28
rect 103 -29 104 -28
rect 104 -29 105 -28
rect 105 -29 106 -28
rect 106 -29 107 -28
rect 107 -29 108 -28
rect 108 -29 109 -28
rect 109 -29 110 -28
rect 110 -29 111 -28
rect 111 -29 112 -28
rect 112 -29 113 -28
rect 113 -29 114 -28
rect 114 -29 115 -28
rect 115 -29 116 -28
rect 116 -29 117 -28
rect 117 -29 118 -28
rect 118 -29 119 -28
rect 119 -29 120 -28
rect 120 -29 121 -28
rect 121 -29 122 -28
rect 122 -29 123 -28
rect 123 -29 124 -28
rect 133 -29 134 -28
rect 134 -29 135 -28
rect 135 -29 136 -28
rect 136 -29 137 -28
rect 137 -29 138 -28
rect 138 -29 139 -28
rect 139 -29 140 -28
rect 140 -29 141 -28
rect 141 -29 142 -28
rect 142 -29 143 -28
rect 143 -29 144 -28
rect 144 -29 145 -28
rect 145 -29 146 -28
rect 146 -29 147 -28
rect 147 -29 148 -28
rect 148 -29 149 -28
rect 149 -29 150 -28
rect 150 -29 151 -28
rect 151 -29 152 -28
rect 152 -29 153 -28
rect 153 -29 154 -28
rect 154 -29 155 -28
rect 155 -29 156 -28
rect 165 -29 166 -28
rect 166 -29 167 -28
rect 167 -29 168 -28
rect 168 -29 169 -28
rect 169 -29 170 -28
rect 170 -29 171 -28
rect 171 -29 172 -28
rect 172 -29 173 -28
rect 173 -29 174 -28
rect 174 -29 175 -28
rect 175 -29 176 -28
rect 176 -29 177 -28
rect 177 -29 178 -28
rect 178 -29 179 -28
rect 179 -29 180 -28
rect 180 -29 181 -28
rect 181 -29 182 -28
rect 182 -29 183 -28
rect 183 -29 184 -28
rect 184 -29 185 -28
rect 185 -29 186 -28
rect 186 -29 187 -28
rect 187 -29 188 -28
rect 188 -29 189 -28
rect 189 -29 190 -28
rect 190 -29 191 -28
rect 191 -29 192 -28
rect 2 -30 3 -29
rect 3 -30 4 -29
rect 4 -30 5 -29
rect 5 -30 6 -29
rect 6 -30 7 -29
rect 7 -30 8 -29
rect 8 -30 9 -29
rect 9 -30 10 -29
rect 10 -30 11 -29
rect 11 -30 12 -29
rect 12 -30 13 -29
rect 13 -30 14 -29
rect 14 -30 15 -29
rect 15 -30 16 -29
rect 16 -30 17 -29
rect 17 -30 18 -29
rect 18 -30 19 -29
rect 19 -30 20 -29
rect 20 -30 21 -29
rect 21 -30 22 -29
rect 22 -30 23 -29
rect 23 -30 24 -29
rect 24 -30 25 -29
rect 25 -30 26 -29
rect 26 -30 27 -29
rect 27 -30 28 -29
rect 37 -30 38 -29
rect 38 -30 39 -29
rect 39 -30 40 -29
rect 40 -30 41 -29
rect 41 -30 42 -29
rect 42 -30 43 -29
rect 43 -30 44 -29
rect 44 -30 45 -29
rect 45 -30 46 -29
rect 46 -30 47 -29
rect 47 -30 48 -29
rect 48 -30 49 -29
rect 49 -30 50 -29
rect 50 -30 51 -29
rect 51 -30 52 -29
rect 52 -30 53 -29
rect 53 -30 54 -29
rect 54 -30 55 -29
rect 55 -30 56 -29
rect 56 -30 57 -29
rect 57 -30 58 -29
rect 58 -30 59 -29
rect 59 -30 60 -29
rect 69 -30 70 -29
rect 70 -30 71 -29
rect 71 -30 72 -29
rect 72 -30 73 -29
rect 73 -30 74 -29
rect 74 -30 75 -29
rect 75 -30 76 -29
rect 76 -30 77 -29
rect 77 -30 78 -29
rect 78 -30 79 -29
rect 79 -30 80 -29
rect 80 -30 81 -29
rect 81 -30 82 -29
rect 82 -30 83 -29
rect 83 -30 84 -29
rect 84 -30 85 -29
rect 85 -30 86 -29
rect 86 -30 87 -29
rect 87 -30 88 -29
rect 88 -30 89 -29
rect 89 -30 90 -29
rect 90 -30 91 -29
rect 91 -30 92 -29
rect 101 -30 102 -29
rect 102 -30 103 -29
rect 103 -30 104 -29
rect 104 -30 105 -29
rect 105 -30 106 -29
rect 106 -30 107 -29
rect 107 -30 108 -29
rect 108 -30 109 -29
rect 109 -30 110 -29
rect 110 -30 111 -29
rect 111 -30 112 -29
rect 112 -30 113 -29
rect 113 -30 114 -29
rect 114 -30 115 -29
rect 115 -30 116 -29
rect 116 -30 117 -29
rect 117 -30 118 -29
rect 118 -30 119 -29
rect 119 -30 120 -29
rect 120 -30 121 -29
rect 121 -30 122 -29
rect 122 -30 123 -29
rect 123 -30 124 -29
rect 133 -30 134 -29
rect 134 -30 135 -29
rect 135 -30 136 -29
rect 136 -30 137 -29
rect 137 -30 138 -29
rect 138 -30 139 -29
rect 139 -30 140 -29
rect 140 -30 141 -29
rect 141 -30 142 -29
rect 142 -30 143 -29
rect 143 -30 144 -29
rect 144 -30 145 -29
rect 145 -30 146 -29
rect 146 -30 147 -29
rect 147 -30 148 -29
rect 148 -30 149 -29
rect 149 -30 150 -29
rect 150 -30 151 -29
rect 151 -30 152 -29
rect 152 -30 153 -29
rect 153 -30 154 -29
rect 154 -30 155 -29
rect 155 -30 156 -29
rect 165 -30 166 -29
rect 166 -30 167 -29
rect 167 -30 168 -29
rect 168 -30 169 -29
rect 169 -30 170 -29
rect 170 -30 171 -29
rect 171 -30 172 -29
rect 172 -30 173 -29
rect 173 -30 174 -29
rect 174 -30 175 -29
rect 175 -30 176 -29
rect 176 -30 177 -29
rect 177 -30 178 -29
rect 178 -30 179 -29
rect 179 -30 180 -29
rect 180 -30 181 -29
rect 181 -30 182 -29
rect 182 -30 183 -29
rect 183 -30 184 -29
rect 184 -30 185 -29
rect 185 -30 186 -29
rect 186 -30 187 -29
rect 187 -30 188 -29
rect 188 -30 189 -29
rect 189 -30 190 -29
rect 190 -30 191 -29
rect 191 -30 192 -29
rect 2 -31 3 -30
rect 3 -31 4 -30
rect 4 -31 5 -30
rect 5 -31 6 -30
rect 6 -31 7 -30
rect 7 -31 8 -30
rect 8 -31 9 -30
rect 9 -31 10 -30
rect 10 -31 11 -30
rect 11 -31 12 -30
rect 12 -31 13 -30
rect 13 -31 14 -30
rect 14 -31 15 -30
rect 15 -31 16 -30
rect 16 -31 17 -30
rect 17 -31 18 -30
rect 18 -31 19 -30
rect 19 -31 20 -30
rect 20 -31 21 -30
rect 21 -31 22 -30
rect 22 -31 23 -30
rect 23 -31 24 -30
rect 24 -31 25 -30
rect 25 -31 26 -30
rect 26 -31 27 -30
rect 27 -31 28 -30
rect 37 -31 38 -30
rect 38 -31 39 -30
rect 39 -31 40 -30
rect 40 -31 41 -30
rect 41 -31 42 -30
rect 42 -31 43 -30
rect 43 -31 44 -30
rect 44 -31 45 -30
rect 45 -31 46 -30
rect 46 -31 47 -30
rect 47 -31 48 -30
rect 48 -31 49 -30
rect 49 -31 50 -30
rect 50 -31 51 -30
rect 51 -31 52 -30
rect 52 -31 53 -30
rect 53 -31 54 -30
rect 54 -31 55 -30
rect 55 -31 56 -30
rect 56 -31 57 -30
rect 57 -31 58 -30
rect 58 -31 59 -30
rect 59 -31 60 -30
rect 69 -31 70 -30
rect 70 -31 71 -30
rect 71 -31 72 -30
rect 72 -31 73 -30
rect 73 -31 74 -30
rect 74 -31 75 -30
rect 75 -31 76 -30
rect 76 -31 77 -30
rect 77 -31 78 -30
rect 78 -31 79 -30
rect 79 -31 80 -30
rect 80 -31 81 -30
rect 81 -31 82 -30
rect 82 -31 83 -30
rect 83 -31 84 -30
rect 84 -31 85 -30
rect 85 -31 86 -30
rect 86 -31 87 -30
rect 87 -31 88 -30
rect 88 -31 89 -30
rect 89 -31 90 -30
rect 90 -31 91 -30
rect 91 -31 92 -30
rect 101 -31 102 -30
rect 102 -31 103 -30
rect 103 -31 104 -30
rect 104 -31 105 -30
rect 105 -31 106 -30
rect 106 -31 107 -30
rect 107 -31 108 -30
rect 108 -31 109 -30
rect 109 -31 110 -30
rect 110 -31 111 -30
rect 111 -31 112 -30
rect 112 -31 113 -30
rect 113 -31 114 -30
rect 114 -31 115 -30
rect 115 -31 116 -30
rect 116 -31 117 -30
rect 117 -31 118 -30
rect 118 -31 119 -30
rect 119 -31 120 -30
rect 120 -31 121 -30
rect 121 -31 122 -30
rect 122 -31 123 -30
rect 123 -31 124 -30
rect 133 -31 134 -30
rect 134 -31 135 -30
rect 135 -31 136 -30
rect 136 -31 137 -30
rect 137 -31 138 -30
rect 138 -31 139 -30
rect 139 -31 140 -30
rect 140 -31 141 -30
rect 141 -31 142 -30
rect 142 -31 143 -30
rect 143 -31 144 -30
rect 144 -31 145 -30
rect 145 -31 146 -30
rect 146 -31 147 -30
rect 147 -31 148 -30
rect 148 -31 149 -30
rect 149 -31 150 -30
rect 150 -31 151 -30
rect 151 -31 152 -30
rect 152 -31 153 -30
rect 153 -31 154 -30
rect 154 -31 155 -30
rect 155 -31 156 -30
rect 165 -31 166 -30
rect 166 -31 167 -30
rect 167 -31 168 -30
rect 168 -31 169 -30
rect 169 -31 170 -30
rect 170 -31 171 -30
rect 171 -31 172 -30
rect 172 -31 173 -30
rect 173 -31 174 -30
rect 174 -31 175 -30
rect 175 -31 176 -30
rect 176 -31 177 -30
rect 177 -31 178 -30
rect 178 -31 179 -30
rect 179 -31 180 -30
rect 180 -31 181 -30
rect 181 -31 182 -30
rect 182 -31 183 -30
rect 183 -31 184 -30
rect 184 -31 185 -30
rect 185 -31 186 -30
rect 186 -31 187 -30
rect 187 -31 188 -30
rect 188 -31 189 -30
rect 189 -31 190 -30
rect 190 -31 191 -30
rect 191 -31 192 -30
rect 2 -32 3 -31
rect 3 -32 4 -31
rect 4 -32 5 -31
rect 5 -32 6 -31
rect 6 -32 7 -31
rect 7 -32 8 -31
rect 8 -32 9 -31
rect 9 -32 10 -31
rect 10 -32 11 -31
rect 11 -32 12 -31
rect 12 -32 13 -31
rect 13 -32 14 -31
rect 14 -32 15 -31
rect 15 -32 16 -31
rect 16 -32 17 -31
rect 17 -32 18 -31
rect 18 -32 19 -31
rect 19 -32 20 -31
rect 20 -32 21 -31
rect 21 -32 22 -31
rect 22 -32 23 -31
rect 23 -32 24 -31
rect 24 -32 25 -31
rect 25 -32 26 -31
rect 26 -32 27 -31
rect 27 -32 28 -31
rect 32 -32 33 -31
rect 33 -32 34 -31
rect 37 -32 38 -31
rect 38 -32 39 -31
rect 39 -32 40 -31
rect 40 -32 41 -31
rect 41 -32 42 -31
rect 42 -32 43 -31
rect 43 -32 44 -31
rect 44 -32 45 -31
rect 45 -32 46 -31
rect 46 -32 47 -31
rect 47 -32 48 -31
rect 48 -32 49 -31
rect 49 -32 50 -31
rect 50 -32 51 -31
rect 51 -32 52 -31
rect 52 -32 53 -31
rect 53 -32 54 -31
rect 54 -32 55 -31
rect 55 -32 56 -31
rect 56 -32 57 -31
rect 57 -32 58 -31
rect 58 -32 59 -31
rect 59 -32 60 -31
rect 64 -32 65 -31
rect 65 -32 66 -31
rect 69 -32 70 -31
rect 70 -32 71 -31
rect 71 -32 72 -31
rect 72 -32 73 -31
rect 73 -32 74 -31
rect 74 -32 75 -31
rect 75 -32 76 -31
rect 76 -32 77 -31
rect 77 -32 78 -31
rect 78 -32 79 -31
rect 79 -32 80 -31
rect 80 -32 81 -31
rect 81 -32 82 -31
rect 82 -32 83 -31
rect 83 -32 84 -31
rect 84 -32 85 -31
rect 85 -32 86 -31
rect 86 -32 87 -31
rect 87 -32 88 -31
rect 88 -32 89 -31
rect 89 -32 90 -31
rect 90 -32 91 -31
rect 91 -32 92 -31
rect 96 -32 97 -31
rect 97 -32 98 -31
rect 101 -32 102 -31
rect 102 -32 103 -31
rect 103 -32 104 -31
rect 104 -32 105 -31
rect 105 -32 106 -31
rect 106 -32 107 -31
rect 107 -32 108 -31
rect 108 -32 109 -31
rect 109 -32 110 -31
rect 110 -32 111 -31
rect 111 -32 112 -31
rect 112 -32 113 -31
rect 113 -32 114 -31
rect 114 -32 115 -31
rect 115 -32 116 -31
rect 116 -32 117 -31
rect 117 -32 118 -31
rect 118 -32 119 -31
rect 119 -32 120 -31
rect 120 -32 121 -31
rect 121 -32 122 -31
rect 122 -32 123 -31
rect 123 -32 124 -31
rect 128 -32 129 -31
rect 129 -32 130 -31
rect 133 -32 134 -31
rect 134 -32 135 -31
rect 135 -32 136 -31
rect 136 -32 137 -31
rect 137 -32 138 -31
rect 138 -32 139 -31
rect 139 -32 140 -31
rect 140 -32 141 -31
rect 141 -32 142 -31
rect 142 -32 143 -31
rect 143 -32 144 -31
rect 144 -32 145 -31
rect 145 -32 146 -31
rect 146 -32 147 -31
rect 147 -32 148 -31
rect 148 -32 149 -31
rect 149 -32 150 -31
rect 150 -32 151 -31
rect 151 -32 152 -31
rect 152 -32 153 -31
rect 153 -32 154 -31
rect 154 -32 155 -31
rect 155 -32 156 -31
rect 160 -32 161 -31
rect 161 -32 162 -31
rect 165 -32 166 -31
rect 166 -32 167 -31
rect 167 -32 168 -31
rect 168 -32 169 -31
rect 169 -32 170 -31
rect 170 -32 171 -31
rect 171 -32 172 -31
rect 172 -32 173 -31
rect 173 -32 174 -31
rect 174 -32 175 -31
rect 175 -32 176 -31
rect 176 -32 177 -31
rect 177 -32 178 -31
rect 178 -32 179 -31
rect 179 -32 180 -31
rect 180 -32 181 -31
rect 181 -32 182 -31
rect 182 -32 183 -31
rect 183 -32 184 -31
rect 184 -32 185 -31
rect 185 -32 186 -31
rect 186 -32 187 -31
rect 187 -32 188 -31
rect 188 -32 189 -31
rect 189 -32 190 -31
rect 190 -32 191 -31
rect 191 -32 192 -31
rect 2 -33 3 -32
rect 3 -33 4 -32
rect 4 -33 5 -32
rect 5 -33 6 -32
rect 6 -33 7 -32
rect 7 -33 8 -32
rect 8 -33 9 -32
rect 9 -33 10 -32
rect 10 -33 11 -32
rect 11 -33 12 -32
rect 12 -33 13 -32
rect 13 -33 14 -32
rect 14 -33 15 -32
rect 18 -33 19 -32
rect 19 -33 20 -32
rect 20 -33 21 -32
rect 21 -33 22 -32
rect 22 -33 23 -32
rect 23 -33 24 -32
rect 24 -33 25 -32
rect 25 -33 26 -32
rect 26 -33 27 -32
rect 27 -33 28 -32
rect 30 -33 31 -32
rect 31 -33 32 -32
rect 32 -33 33 -32
rect 33 -33 34 -32
rect 34 -33 35 -32
rect 37 -33 38 -32
rect 38 -33 39 -32
rect 39 -33 40 -32
rect 40 -33 41 -32
rect 41 -33 42 -32
rect 42 -33 43 -32
rect 43 -33 44 -32
rect 44 -33 45 -32
rect 45 -33 46 -32
rect 46 -33 47 -32
rect 50 -33 51 -32
rect 51 -33 52 -32
rect 52 -33 53 -32
rect 53 -33 54 -32
rect 54 -33 55 -32
rect 55 -33 56 -32
rect 56 -33 57 -32
rect 57 -33 58 -32
rect 58 -33 59 -32
rect 59 -33 60 -32
rect 62 -33 63 -32
rect 63 -33 64 -32
rect 64 -33 65 -32
rect 65 -33 66 -32
rect 66 -33 67 -32
rect 69 -33 70 -32
rect 70 -33 71 -32
rect 71 -33 72 -32
rect 72 -33 73 -32
rect 73 -33 74 -32
rect 74 -33 75 -32
rect 75 -33 76 -32
rect 76 -33 77 -32
rect 77 -33 78 -32
rect 78 -33 79 -32
rect 82 -33 83 -32
rect 83 -33 84 -32
rect 84 -33 85 -32
rect 85 -33 86 -32
rect 86 -33 87 -32
rect 87 -33 88 -32
rect 88 -33 89 -32
rect 89 -33 90 -32
rect 90 -33 91 -32
rect 91 -33 92 -32
rect 94 -33 95 -32
rect 95 -33 96 -32
rect 96 -33 97 -32
rect 97 -33 98 -32
rect 98 -33 99 -32
rect 101 -33 102 -32
rect 102 -33 103 -32
rect 103 -33 104 -32
rect 104 -33 105 -32
rect 105 -33 106 -32
rect 106 -33 107 -32
rect 107 -33 108 -32
rect 108 -33 109 -32
rect 109 -33 110 -32
rect 110 -33 111 -32
rect 114 -33 115 -32
rect 115 -33 116 -32
rect 116 -33 117 -32
rect 117 -33 118 -32
rect 118 -33 119 -32
rect 119 -33 120 -32
rect 120 -33 121 -32
rect 121 -33 122 -32
rect 122 -33 123 -32
rect 123 -33 124 -32
rect 126 -33 127 -32
rect 127 -33 128 -32
rect 128 -33 129 -32
rect 129 -33 130 -32
rect 130 -33 131 -32
rect 133 -33 134 -32
rect 134 -33 135 -32
rect 135 -33 136 -32
rect 136 -33 137 -32
rect 137 -33 138 -32
rect 138 -33 139 -32
rect 139 -33 140 -32
rect 140 -33 141 -32
rect 141 -33 142 -32
rect 142 -33 143 -32
rect 146 -33 147 -32
rect 147 -33 148 -32
rect 148 -33 149 -32
rect 149 -33 150 -32
rect 150 -33 151 -32
rect 151 -33 152 -32
rect 152 -33 153 -32
rect 153 -33 154 -32
rect 154 -33 155 -32
rect 155 -33 156 -32
rect 158 -33 159 -32
rect 159 -33 160 -32
rect 160 -33 161 -32
rect 161 -33 162 -32
rect 162 -33 163 -32
rect 165 -33 166 -32
rect 166 -33 167 -32
rect 167 -33 168 -32
rect 168 -33 169 -32
rect 169 -33 170 -32
rect 170 -33 171 -32
rect 171 -33 172 -32
rect 172 -33 173 -32
rect 173 -33 174 -32
rect 174 -33 175 -32
rect 178 -33 179 -32
rect 179 -33 180 -32
rect 180 -33 181 -32
rect 181 -33 182 -32
rect 182 -33 183 -32
rect 183 -33 184 -32
rect 184 -33 185 -32
rect 185 -33 186 -32
rect 186 -33 187 -32
rect 187 -33 188 -32
rect 188 -33 189 -32
rect 189 -33 190 -32
rect 190 -33 191 -32
rect 191 -33 192 -32
rect 2 -34 3 -33
rect 3 -34 4 -33
rect 4 -34 5 -33
rect 5 -34 6 -33
rect 6 -34 7 -33
rect 7 -34 8 -33
rect 8 -34 9 -33
rect 9 -34 10 -33
rect 10 -34 11 -33
rect 11 -34 12 -33
rect 12 -34 13 -33
rect 13 -34 14 -33
rect 14 -34 15 -33
rect 18 -34 19 -33
rect 19 -34 20 -33
rect 20 -34 21 -33
rect 21 -34 22 -33
rect 22 -34 23 -33
rect 23 -34 24 -33
rect 24 -34 25 -33
rect 25 -34 26 -33
rect 26 -34 27 -33
rect 27 -34 28 -33
rect 28 -34 29 -33
rect 29 -34 30 -33
rect 30 -34 31 -33
rect 31 -34 32 -33
rect 32 -34 33 -33
rect 33 -34 34 -33
rect 34 -34 35 -33
rect 35 -34 36 -33
rect 36 -34 37 -33
rect 37 -34 38 -33
rect 38 -34 39 -33
rect 39 -34 40 -33
rect 40 -34 41 -33
rect 41 -34 42 -33
rect 42 -34 43 -33
rect 43 -34 44 -33
rect 44 -34 45 -33
rect 45 -34 46 -33
rect 46 -34 47 -33
rect 50 -34 51 -33
rect 51 -34 52 -33
rect 52 -34 53 -33
rect 53 -34 54 -33
rect 54 -34 55 -33
rect 55 -34 56 -33
rect 56 -34 57 -33
rect 57 -34 58 -33
rect 58 -34 59 -33
rect 59 -34 60 -33
rect 60 -34 61 -33
rect 61 -34 62 -33
rect 62 -34 63 -33
rect 63 -34 64 -33
rect 64 -34 65 -33
rect 65 -34 66 -33
rect 66 -34 67 -33
rect 67 -34 68 -33
rect 68 -34 69 -33
rect 69 -34 70 -33
rect 70 -34 71 -33
rect 71 -34 72 -33
rect 72 -34 73 -33
rect 73 -34 74 -33
rect 74 -34 75 -33
rect 75 -34 76 -33
rect 76 -34 77 -33
rect 77 -34 78 -33
rect 78 -34 79 -33
rect 82 -34 83 -33
rect 83 -34 84 -33
rect 84 -34 85 -33
rect 85 -34 86 -33
rect 86 -34 87 -33
rect 87 -34 88 -33
rect 88 -34 89 -33
rect 89 -34 90 -33
rect 90 -34 91 -33
rect 91 -34 92 -33
rect 92 -34 93 -33
rect 93 -34 94 -33
rect 94 -34 95 -33
rect 95 -34 96 -33
rect 96 -34 97 -33
rect 97 -34 98 -33
rect 98 -34 99 -33
rect 99 -34 100 -33
rect 100 -34 101 -33
rect 101 -34 102 -33
rect 102 -34 103 -33
rect 103 -34 104 -33
rect 104 -34 105 -33
rect 105 -34 106 -33
rect 106 -34 107 -33
rect 107 -34 108 -33
rect 108 -34 109 -33
rect 109 -34 110 -33
rect 110 -34 111 -33
rect 114 -34 115 -33
rect 115 -34 116 -33
rect 116 -34 117 -33
rect 117 -34 118 -33
rect 118 -34 119 -33
rect 119 -34 120 -33
rect 120 -34 121 -33
rect 121 -34 122 -33
rect 122 -34 123 -33
rect 123 -34 124 -33
rect 124 -34 125 -33
rect 125 -34 126 -33
rect 126 -34 127 -33
rect 127 -34 128 -33
rect 128 -34 129 -33
rect 129 -34 130 -33
rect 130 -34 131 -33
rect 131 -34 132 -33
rect 132 -34 133 -33
rect 133 -34 134 -33
rect 134 -34 135 -33
rect 135 -34 136 -33
rect 136 -34 137 -33
rect 137 -34 138 -33
rect 138 -34 139 -33
rect 139 -34 140 -33
rect 140 -34 141 -33
rect 141 -34 142 -33
rect 142 -34 143 -33
rect 146 -34 147 -33
rect 147 -34 148 -33
rect 148 -34 149 -33
rect 149 -34 150 -33
rect 150 -34 151 -33
rect 151 -34 152 -33
rect 152 -34 153 -33
rect 153 -34 154 -33
rect 154 -34 155 -33
rect 155 -34 156 -33
rect 156 -34 157 -33
rect 157 -34 158 -33
rect 158 -34 159 -33
rect 159 -34 160 -33
rect 160 -34 161 -33
rect 161 -34 162 -33
rect 162 -34 163 -33
rect 163 -34 164 -33
rect 164 -34 165 -33
rect 165 -34 166 -33
rect 166 -34 167 -33
rect 167 -34 168 -33
rect 168 -34 169 -33
rect 169 -34 170 -33
rect 170 -34 171 -33
rect 171 -34 172 -33
rect 172 -34 173 -33
rect 173 -34 174 -33
rect 174 -34 175 -33
rect 178 -34 179 -33
rect 179 -34 180 -33
rect 180 -34 181 -33
rect 181 -34 182 -33
rect 182 -34 183 -33
rect 183 -34 184 -33
rect 184 -34 185 -33
rect 185 -34 186 -33
rect 186 -34 187 -33
rect 187 -34 188 -33
rect 188 -34 189 -33
rect 189 -34 190 -33
rect 190 -34 191 -33
rect 191 -34 192 -33
rect 2 -35 3 -34
rect 3 -35 4 -34
rect 4 -35 5 -34
rect 5 -35 6 -34
rect 6 -35 7 -34
rect 7 -35 8 -34
rect 8 -35 9 -34
rect 9 -35 10 -34
rect 10 -35 11 -34
rect 11 -35 12 -34
rect 12 -35 13 -34
rect 13 -35 14 -34
rect 14 -35 15 -34
rect 19 -35 20 -34
rect 20 -35 21 -34
rect 21 -35 22 -34
rect 22 -35 23 -34
rect 23 -35 24 -34
rect 24 -35 25 -34
rect 25 -35 26 -34
rect 26 -35 27 -34
rect 27 -35 28 -34
rect 28 -35 29 -34
rect 29 -35 30 -34
rect 30 -35 31 -34
rect 31 -35 32 -34
rect 32 -35 33 -34
rect 33 -35 34 -34
rect 34 -35 35 -34
rect 35 -35 36 -34
rect 36 -35 37 -34
rect 37 -35 38 -34
rect 38 -35 39 -34
rect 39 -35 40 -34
rect 40 -35 41 -34
rect 41 -35 42 -34
rect 42 -35 43 -34
rect 43 -35 44 -34
rect 44 -35 45 -34
rect 45 -35 46 -34
rect 46 -35 47 -34
rect 51 -35 52 -34
rect 52 -35 53 -34
rect 53 -35 54 -34
rect 54 -35 55 -34
rect 55 -35 56 -34
rect 56 -35 57 -34
rect 57 -35 58 -34
rect 58 -35 59 -34
rect 59 -35 60 -34
rect 60 -35 61 -34
rect 61 -35 62 -34
rect 62 -35 63 -34
rect 63 -35 64 -34
rect 64 -35 65 -34
rect 65 -35 66 -34
rect 66 -35 67 -34
rect 67 -35 68 -34
rect 68 -35 69 -34
rect 69 -35 70 -34
rect 70 -35 71 -34
rect 71 -35 72 -34
rect 72 -35 73 -34
rect 73 -35 74 -34
rect 74 -35 75 -34
rect 75 -35 76 -34
rect 76 -35 77 -34
rect 77 -35 78 -34
rect 78 -35 79 -34
rect 83 -35 84 -34
rect 84 -35 85 -34
rect 85 -35 86 -34
rect 86 -35 87 -34
rect 87 -35 88 -34
rect 88 -35 89 -34
rect 89 -35 90 -34
rect 90 -35 91 -34
rect 91 -35 92 -34
rect 92 -35 93 -34
rect 93 -35 94 -34
rect 94 -35 95 -34
rect 95 -35 96 -34
rect 96 -35 97 -34
rect 97 -35 98 -34
rect 98 -35 99 -34
rect 99 -35 100 -34
rect 100 -35 101 -34
rect 101 -35 102 -34
rect 102 -35 103 -34
rect 103 -35 104 -34
rect 104 -35 105 -34
rect 105 -35 106 -34
rect 106 -35 107 -34
rect 107 -35 108 -34
rect 108 -35 109 -34
rect 109 -35 110 -34
rect 110 -35 111 -34
rect 115 -35 116 -34
rect 116 -35 117 -34
rect 117 -35 118 -34
rect 118 -35 119 -34
rect 119 -35 120 -34
rect 120 -35 121 -34
rect 121 -35 122 -34
rect 122 -35 123 -34
rect 123 -35 124 -34
rect 124 -35 125 -34
rect 125 -35 126 -34
rect 126 -35 127 -34
rect 127 -35 128 -34
rect 128 -35 129 -34
rect 129 -35 130 -34
rect 130 -35 131 -34
rect 131 -35 132 -34
rect 132 -35 133 -34
rect 133 -35 134 -34
rect 134 -35 135 -34
rect 135 -35 136 -34
rect 136 -35 137 -34
rect 137 -35 138 -34
rect 138 -35 139 -34
rect 139 -35 140 -34
rect 140 -35 141 -34
rect 141 -35 142 -34
rect 142 -35 143 -34
rect 147 -35 148 -34
rect 148 -35 149 -34
rect 149 -35 150 -34
rect 150 -35 151 -34
rect 151 -35 152 -34
rect 152 -35 153 -34
rect 153 -35 154 -34
rect 154 -35 155 -34
rect 155 -35 156 -34
rect 156 -35 157 -34
rect 157 -35 158 -34
rect 158 -35 159 -34
rect 159 -35 160 -34
rect 160 -35 161 -34
rect 161 -35 162 -34
rect 162 -35 163 -34
rect 163 -35 164 -34
rect 164 -35 165 -34
rect 165 -35 166 -34
rect 166 -35 167 -34
rect 167 -35 168 -34
rect 168 -35 169 -34
rect 169 -35 170 -34
rect 170 -35 171 -34
rect 171 -35 172 -34
rect 172 -35 173 -34
rect 173 -35 174 -34
rect 174 -35 175 -34
rect 179 -35 180 -34
rect 180 -35 181 -34
rect 181 -35 182 -34
rect 182 -35 183 -34
rect 183 -35 184 -34
rect 184 -35 185 -34
rect 185 -35 186 -34
rect 186 -35 187 -34
rect 187 -35 188 -34
rect 188 -35 189 -34
rect 189 -35 190 -34
rect 190 -35 191 -34
rect 191 -35 192 -34
rect 2 -36 3 -35
rect 3 -36 4 -35
rect 4 -36 5 -35
rect 5 -36 6 -35
rect 6 -36 7 -35
rect 7 -36 8 -35
rect 8 -36 9 -35
rect 9 -36 10 -35
rect 10 -36 11 -35
rect 11 -36 12 -35
rect 12 -36 13 -35
rect 13 -36 14 -35
rect 14 -36 15 -35
rect 19 -36 20 -35
rect 20 -36 21 -35
rect 21 -36 22 -35
rect 22 -36 23 -35
rect 23 -36 24 -35
rect 24 -36 25 -35
rect 25 -36 26 -35
rect 26 -36 27 -35
rect 27 -36 28 -35
rect 28 -36 29 -35
rect 29 -36 30 -35
rect 30 -36 31 -35
rect 31 -36 32 -35
rect 32 -36 33 -35
rect 33 -36 34 -35
rect 34 -36 35 -35
rect 35 -36 36 -35
rect 36 -36 37 -35
rect 37 -36 38 -35
rect 38 -36 39 -35
rect 39 -36 40 -35
rect 40 -36 41 -35
rect 41 -36 42 -35
rect 42 -36 43 -35
rect 43 -36 44 -35
rect 44 -36 45 -35
rect 45 -36 46 -35
rect 46 -36 47 -35
rect 51 -36 52 -35
rect 52 -36 53 -35
rect 53 -36 54 -35
rect 54 -36 55 -35
rect 55 -36 56 -35
rect 56 -36 57 -35
rect 57 -36 58 -35
rect 58 -36 59 -35
rect 59 -36 60 -35
rect 60 -36 61 -35
rect 61 -36 62 -35
rect 62 -36 63 -35
rect 63 -36 64 -35
rect 64 -36 65 -35
rect 65 -36 66 -35
rect 66 -36 67 -35
rect 67 -36 68 -35
rect 68 -36 69 -35
rect 69 -36 70 -35
rect 70 -36 71 -35
rect 71 -36 72 -35
rect 72 -36 73 -35
rect 73 -36 74 -35
rect 74 -36 75 -35
rect 75 -36 76 -35
rect 76 -36 77 -35
rect 77 -36 78 -35
rect 78 -36 79 -35
rect 83 -36 84 -35
rect 84 -36 85 -35
rect 85 -36 86 -35
rect 86 -36 87 -35
rect 87 -36 88 -35
rect 88 -36 89 -35
rect 89 -36 90 -35
rect 90 -36 91 -35
rect 91 -36 92 -35
rect 92 -36 93 -35
rect 93 -36 94 -35
rect 94 -36 95 -35
rect 95 -36 96 -35
rect 96 -36 97 -35
rect 97 -36 98 -35
rect 98 -36 99 -35
rect 99 -36 100 -35
rect 100 -36 101 -35
rect 101 -36 102 -35
rect 102 -36 103 -35
rect 103 -36 104 -35
rect 104 -36 105 -35
rect 105 -36 106 -35
rect 106 -36 107 -35
rect 107 -36 108 -35
rect 108 -36 109 -35
rect 109 -36 110 -35
rect 110 -36 111 -35
rect 115 -36 116 -35
rect 116 -36 117 -35
rect 117 -36 118 -35
rect 118 -36 119 -35
rect 119 -36 120 -35
rect 120 -36 121 -35
rect 121 -36 122 -35
rect 122 -36 123 -35
rect 123 -36 124 -35
rect 124 -36 125 -35
rect 125 -36 126 -35
rect 126 -36 127 -35
rect 127 -36 128 -35
rect 128 -36 129 -35
rect 129 -36 130 -35
rect 130 -36 131 -35
rect 131 -36 132 -35
rect 132 -36 133 -35
rect 133 -36 134 -35
rect 134 -36 135 -35
rect 135 -36 136 -35
rect 136 -36 137 -35
rect 137 -36 138 -35
rect 138 -36 139 -35
rect 139 -36 140 -35
rect 140 -36 141 -35
rect 141 -36 142 -35
rect 142 -36 143 -35
rect 147 -36 148 -35
rect 148 -36 149 -35
rect 149 -36 150 -35
rect 150 -36 151 -35
rect 151 -36 152 -35
rect 152 -36 153 -35
rect 153 -36 154 -35
rect 154 -36 155 -35
rect 155 -36 156 -35
rect 156 -36 157 -35
rect 157 -36 158 -35
rect 158 -36 159 -35
rect 159 -36 160 -35
rect 160 -36 161 -35
rect 161 -36 162 -35
rect 162 -36 163 -35
rect 163 -36 164 -35
rect 164 -36 165 -35
rect 165 -36 166 -35
rect 166 -36 167 -35
rect 167 -36 168 -35
rect 168 -36 169 -35
rect 169 -36 170 -35
rect 170 -36 171 -35
rect 171 -36 172 -35
rect 172 -36 173 -35
rect 173 -36 174 -35
rect 174 -36 175 -35
rect 179 -36 180 -35
rect 180 -36 181 -35
rect 181 -36 182 -35
rect 182 -36 183 -35
rect 183 -36 184 -35
rect 184 -36 185 -35
rect 185 -36 186 -35
rect 186 -36 187 -35
rect 187 -36 188 -35
rect 188 -36 189 -35
rect 189 -36 190 -35
rect 190 -36 191 -35
rect 191 -36 192 -35
rect 2 -37 3 -36
rect 3 -37 4 -36
rect 4 -37 5 -36
rect 5 -37 6 -36
rect 6 -37 7 -36
rect 7 -37 8 -36
rect 8 -37 9 -36
rect 9 -37 10 -36
rect 10 -37 11 -36
rect 11 -37 12 -36
rect 12 -37 13 -36
rect 13 -37 14 -36
rect 19 -37 20 -36
rect 20 -37 21 -36
rect 21 -37 22 -36
rect 22 -37 23 -36
rect 23 -37 24 -36
rect 24 -37 25 -36
rect 25 -37 26 -36
rect 26 -37 27 -36
rect 27 -37 28 -36
rect 28 -37 29 -36
rect 29 -37 30 -36
rect 30 -37 31 -36
rect 31 -37 32 -36
rect 32 -37 33 -36
rect 33 -37 34 -36
rect 34 -37 35 -36
rect 35 -37 36 -36
rect 36 -37 37 -36
rect 37 -37 38 -36
rect 38 -37 39 -36
rect 39 -37 40 -36
rect 40 -37 41 -36
rect 41 -37 42 -36
rect 42 -37 43 -36
rect 43 -37 44 -36
rect 44 -37 45 -36
rect 45 -37 46 -36
rect 51 -37 52 -36
rect 52 -37 53 -36
rect 53 -37 54 -36
rect 54 -37 55 -36
rect 55 -37 56 -36
rect 56 -37 57 -36
rect 57 -37 58 -36
rect 58 -37 59 -36
rect 59 -37 60 -36
rect 60 -37 61 -36
rect 61 -37 62 -36
rect 62 -37 63 -36
rect 63 -37 64 -36
rect 64 -37 65 -36
rect 65 -37 66 -36
rect 66 -37 67 -36
rect 67 -37 68 -36
rect 68 -37 69 -36
rect 69 -37 70 -36
rect 70 -37 71 -36
rect 71 -37 72 -36
rect 72 -37 73 -36
rect 73 -37 74 -36
rect 74 -37 75 -36
rect 75 -37 76 -36
rect 76 -37 77 -36
rect 77 -37 78 -36
rect 83 -37 84 -36
rect 84 -37 85 -36
rect 85 -37 86 -36
rect 86 -37 87 -36
rect 87 -37 88 -36
rect 88 -37 89 -36
rect 89 -37 90 -36
rect 90 -37 91 -36
rect 91 -37 92 -36
rect 92 -37 93 -36
rect 93 -37 94 -36
rect 94 -37 95 -36
rect 95 -37 96 -36
rect 96 -37 97 -36
rect 97 -37 98 -36
rect 98 -37 99 -36
rect 99 -37 100 -36
rect 100 -37 101 -36
rect 101 -37 102 -36
rect 102 -37 103 -36
rect 103 -37 104 -36
rect 104 -37 105 -36
rect 105 -37 106 -36
rect 106 -37 107 -36
rect 107 -37 108 -36
rect 108 -37 109 -36
rect 109 -37 110 -36
rect 115 -37 116 -36
rect 116 -37 117 -36
rect 117 -37 118 -36
rect 118 -37 119 -36
rect 119 -37 120 -36
rect 120 -37 121 -36
rect 121 -37 122 -36
rect 122 -37 123 -36
rect 123 -37 124 -36
rect 124 -37 125 -36
rect 125 -37 126 -36
rect 126 -37 127 -36
rect 127 -37 128 -36
rect 128 -37 129 -36
rect 129 -37 130 -36
rect 130 -37 131 -36
rect 131 -37 132 -36
rect 132 -37 133 -36
rect 133 -37 134 -36
rect 134 -37 135 -36
rect 135 -37 136 -36
rect 136 -37 137 -36
rect 137 -37 138 -36
rect 138 -37 139 -36
rect 139 -37 140 -36
rect 140 -37 141 -36
rect 141 -37 142 -36
rect 147 -37 148 -36
rect 148 -37 149 -36
rect 149 -37 150 -36
rect 150 -37 151 -36
rect 151 -37 152 -36
rect 152 -37 153 -36
rect 153 -37 154 -36
rect 154 -37 155 -36
rect 155 -37 156 -36
rect 156 -37 157 -36
rect 157 -37 158 -36
rect 158 -37 159 -36
rect 159 -37 160 -36
rect 160 -37 161 -36
rect 161 -37 162 -36
rect 162 -37 163 -36
rect 163 -37 164 -36
rect 164 -37 165 -36
rect 165 -37 166 -36
rect 166 -37 167 -36
rect 167 -37 168 -36
rect 168 -37 169 -36
rect 169 -37 170 -36
rect 170 -37 171 -36
rect 171 -37 172 -36
rect 172 -37 173 -36
rect 173 -37 174 -36
rect 179 -37 180 -36
rect 180 -37 181 -36
rect 181 -37 182 -36
rect 182 -37 183 -36
rect 183 -37 184 -36
rect 184 -37 185 -36
rect 185 -37 186 -36
rect 186 -37 187 -36
rect 187 -37 188 -36
rect 188 -37 189 -36
rect 189 -37 190 -36
rect 190 -37 191 -36
rect 191 -37 192 -36
rect 2 -38 3 -37
rect 3 -38 4 -37
rect 4 -38 5 -37
rect 5 -38 6 -37
rect 6 -38 7 -37
rect 7 -38 8 -37
rect 8 -38 9 -37
rect 25 -38 26 -37
rect 26 -38 27 -37
rect 27 -38 28 -37
rect 28 -38 29 -37
rect 29 -38 30 -37
rect 30 -38 31 -37
rect 31 -38 32 -37
rect 32 -38 33 -37
rect 33 -38 34 -37
rect 34 -38 35 -37
rect 35 -38 36 -37
rect 36 -38 37 -37
rect 37 -38 38 -37
rect 38 -38 39 -37
rect 39 -38 40 -37
rect 40 -38 41 -37
rect 57 -38 58 -37
rect 58 -38 59 -37
rect 59 -38 60 -37
rect 60 -38 61 -37
rect 61 -38 62 -37
rect 62 -38 63 -37
rect 63 -38 64 -37
rect 64 -38 65 -37
rect 65 -38 66 -37
rect 66 -38 67 -37
rect 67 -38 68 -37
rect 68 -38 69 -37
rect 69 -38 70 -37
rect 70 -38 71 -37
rect 71 -38 72 -37
rect 72 -38 73 -37
rect 89 -38 90 -37
rect 90 -38 91 -37
rect 91 -38 92 -37
rect 92 -38 93 -37
rect 93 -38 94 -37
rect 94 -38 95 -37
rect 95 -38 96 -37
rect 96 -38 97 -37
rect 97 -38 98 -37
rect 98 -38 99 -37
rect 99 -38 100 -37
rect 100 -38 101 -37
rect 101 -38 102 -37
rect 102 -38 103 -37
rect 103 -38 104 -37
rect 104 -38 105 -37
rect 121 -38 122 -37
rect 122 -38 123 -37
rect 123 -38 124 -37
rect 124 -38 125 -37
rect 125 -38 126 -37
rect 126 -38 127 -37
rect 127 -38 128 -37
rect 128 -38 129 -37
rect 129 -38 130 -37
rect 130 -38 131 -37
rect 131 -38 132 -37
rect 132 -38 133 -37
rect 133 -38 134 -37
rect 134 -38 135 -37
rect 135 -38 136 -37
rect 136 -38 137 -37
rect 153 -38 154 -37
rect 154 -38 155 -37
rect 155 -38 156 -37
rect 156 -38 157 -37
rect 157 -38 158 -37
rect 158 -38 159 -37
rect 159 -38 160 -37
rect 160 -38 161 -37
rect 161 -38 162 -37
rect 162 -38 163 -37
rect 163 -38 164 -37
rect 164 -38 165 -37
rect 165 -38 166 -37
rect 166 -38 167 -37
rect 167 -38 168 -37
rect 168 -38 169 -37
rect 185 -38 186 -37
rect 186 -38 187 -37
rect 187 -38 188 -37
rect 188 -38 189 -37
rect 189 -38 190 -37
rect 190 -38 191 -37
rect 191 -38 192 -37
rect 2 -39 3 -38
rect 3 -39 4 -38
rect 4 -39 5 -38
rect 5 -39 6 -38
rect 6 -39 7 -38
rect 7 -39 8 -38
rect 8 -39 9 -38
rect 24 -39 25 -38
rect 25 -39 26 -38
rect 26 -39 27 -38
rect 27 -39 28 -38
rect 28 -39 29 -38
rect 29 -39 30 -38
rect 30 -39 31 -38
rect 31 -39 32 -38
rect 32 -39 33 -38
rect 33 -39 34 -38
rect 34 -39 35 -38
rect 35 -39 36 -38
rect 36 -39 37 -38
rect 37 -39 38 -38
rect 38 -39 39 -38
rect 39 -39 40 -38
rect 40 -39 41 -38
rect 56 -39 57 -38
rect 57 -39 58 -38
rect 58 -39 59 -38
rect 59 -39 60 -38
rect 60 -39 61 -38
rect 61 -39 62 -38
rect 62 -39 63 -38
rect 63 -39 64 -38
rect 64 -39 65 -38
rect 65 -39 66 -38
rect 66 -39 67 -38
rect 67 -39 68 -38
rect 68 -39 69 -38
rect 69 -39 70 -38
rect 70 -39 71 -38
rect 71 -39 72 -38
rect 72 -39 73 -38
rect 88 -39 89 -38
rect 89 -39 90 -38
rect 90 -39 91 -38
rect 91 -39 92 -38
rect 92 -39 93 -38
rect 93 -39 94 -38
rect 94 -39 95 -38
rect 95 -39 96 -38
rect 96 -39 97 -38
rect 97 -39 98 -38
rect 98 -39 99 -38
rect 99 -39 100 -38
rect 100 -39 101 -38
rect 101 -39 102 -38
rect 102 -39 103 -38
rect 103 -39 104 -38
rect 104 -39 105 -38
rect 120 -39 121 -38
rect 121 -39 122 -38
rect 122 -39 123 -38
rect 123 -39 124 -38
rect 124 -39 125 -38
rect 125 -39 126 -38
rect 126 -39 127 -38
rect 127 -39 128 -38
rect 128 -39 129 -38
rect 129 -39 130 -38
rect 130 -39 131 -38
rect 131 -39 132 -38
rect 132 -39 133 -38
rect 133 -39 134 -38
rect 134 -39 135 -38
rect 135 -39 136 -38
rect 136 -39 137 -38
rect 152 -39 153 -38
rect 153 -39 154 -38
rect 154 -39 155 -38
rect 155 -39 156 -38
rect 156 -39 157 -38
rect 157 -39 158 -38
rect 158 -39 159 -38
rect 159 -39 160 -38
rect 160 -39 161 -38
rect 161 -39 162 -38
rect 162 -39 163 -38
rect 163 -39 164 -38
rect 164 -39 165 -38
rect 165 -39 166 -38
rect 166 -39 167 -38
rect 167 -39 168 -38
rect 168 -39 169 -38
rect 184 -39 185 -38
rect 185 -39 186 -38
rect 186 -39 187 -38
rect 187 -39 188 -38
rect 188 -39 189 -38
rect 189 -39 190 -38
rect 190 -39 191 -38
rect 191 -39 192 -38
rect 2 -40 3 -39
rect 3 -40 4 -39
rect 4 -40 5 -39
rect 5 -40 6 -39
rect 6 -40 7 -39
rect 7 -40 8 -39
rect 8 -40 9 -39
rect 9 -40 10 -39
rect 23 -40 24 -39
rect 24 -40 25 -39
rect 25 -40 26 -39
rect 26 -40 27 -39
rect 27 -40 28 -39
rect 28 -40 29 -39
rect 29 -40 30 -39
rect 30 -40 31 -39
rect 31 -40 32 -39
rect 32 -40 33 -39
rect 33 -40 34 -39
rect 34 -40 35 -39
rect 35 -40 36 -39
rect 36 -40 37 -39
rect 37 -40 38 -39
rect 38 -40 39 -39
rect 39 -40 40 -39
rect 40 -40 41 -39
rect 41 -40 42 -39
rect 55 -40 56 -39
rect 56 -40 57 -39
rect 57 -40 58 -39
rect 58 -40 59 -39
rect 59 -40 60 -39
rect 60 -40 61 -39
rect 61 -40 62 -39
rect 62 -40 63 -39
rect 63 -40 64 -39
rect 64 -40 65 -39
rect 65 -40 66 -39
rect 66 -40 67 -39
rect 67 -40 68 -39
rect 68 -40 69 -39
rect 69 -40 70 -39
rect 70 -40 71 -39
rect 71 -40 72 -39
rect 72 -40 73 -39
rect 73 -40 74 -39
rect 87 -40 88 -39
rect 88 -40 89 -39
rect 89 -40 90 -39
rect 90 -40 91 -39
rect 91 -40 92 -39
rect 92 -40 93 -39
rect 93 -40 94 -39
rect 94 -40 95 -39
rect 95 -40 96 -39
rect 96 -40 97 -39
rect 97 -40 98 -39
rect 98 -40 99 -39
rect 99 -40 100 -39
rect 100 -40 101 -39
rect 101 -40 102 -39
rect 102 -40 103 -39
rect 103 -40 104 -39
rect 104 -40 105 -39
rect 105 -40 106 -39
rect 119 -40 120 -39
rect 120 -40 121 -39
rect 121 -40 122 -39
rect 122 -40 123 -39
rect 123 -40 124 -39
rect 124 -40 125 -39
rect 125 -40 126 -39
rect 126 -40 127 -39
rect 127 -40 128 -39
rect 128 -40 129 -39
rect 129 -40 130 -39
rect 130 -40 131 -39
rect 131 -40 132 -39
rect 132 -40 133 -39
rect 133 -40 134 -39
rect 134 -40 135 -39
rect 135 -40 136 -39
rect 136 -40 137 -39
rect 137 -40 138 -39
rect 151 -40 152 -39
rect 152 -40 153 -39
rect 153 -40 154 -39
rect 154 -40 155 -39
rect 155 -40 156 -39
rect 156 -40 157 -39
rect 157 -40 158 -39
rect 158 -40 159 -39
rect 159 -40 160 -39
rect 160 -40 161 -39
rect 161 -40 162 -39
rect 162 -40 163 -39
rect 163 -40 164 -39
rect 164 -40 165 -39
rect 165 -40 166 -39
rect 166 -40 167 -39
rect 167 -40 168 -39
rect 168 -40 169 -39
rect 169 -40 170 -39
rect 183 -40 184 -39
rect 184 -40 185 -39
rect 185 -40 186 -39
rect 186 -40 187 -39
rect 187 -40 188 -39
rect 188 -40 189 -39
rect 189 -40 190 -39
rect 190 -40 191 -39
rect 191 -40 192 -39
rect 192 -40 193 -39
rect 193 -40 194 -39
rect 194 -40 195 -39
rect 195 -40 196 -39
rect 196 -40 197 -39
rect 197 -40 198 -39
rect 198 -40 199 -39
rect 199 -40 200 -39
rect 200 -40 201 -39
rect 201 -40 202 -39
rect 202 -40 203 -39
rect 203 -40 204 -39
rect 204 -40 205 -39
rect 205 -40 206 -39
rect 206 -40 207 -39
rect 207 -40 208 -39
rect 208 -40 209 -39
rect 209 -40 210 -39
rect 210 -40 211 -39
rect 211 -40 212 -39
rect 212 -40 213 -39
rect 213 -40 214 -39
rect 214 -40 215 -39
rect 215 -40 216 -39
rect 216 -40 217 -39
rect 217 -40 218 -39
rect 218 -40 219 -39
rect 219 -40 220 -39
rect 220 -40 221 -39
rect 221 -40 222 -39
rect 222 -40 223 -39
rect 223 -40 224 -39
rect 224 -40 225 -39
rect 225 -40 226 -39
rect 226 -40 227 -39
rect 227 -40 228 -39
rect 228 -40 229 -39
rect 229 -40 230 -39
rect 230 -40 231 -39
rect 231 -40 232 -39
rect 232 -40 233 -39
rect 233 -40 234 -39
rect 234 -40 235 -39
rect 235 -40 236 -39
rect 236 -40 237 -39
rect 237 -40 238 -39
rect 238 -40 239 -39
rect 239 -40 240 -39
rect 240 -40 241 -39
rect 241 -40 242 -39
rect 242 -40 243 -39
rect 243 -40 244 -39
rect 244 -40 245 -39
rect 245 -40 246 -39
rect 246 -40 247 -39
rect 247 -40 248 -39
rect 248 -40 249 -39
rect 249 -40 250 -39
rect 250 -40 251 -39
rect 251 -40 252 -39
rect 252 -40 253 -39
rect 253 -40 254 -39
rect 254 -40 255 -39
rect 255 -40 256 -39
rect 256 -40 257 -39
rect 257 -40 258 -39
rect 258 -40 259 -39
rect 259 -40 260 -39
rect 260 -40 261 -39
rect 261 -40 262 -39
rect 262 -40 263 -39
rect 263 -40 264 -39
rect 264 -40 265 -39
rect 265 -40 266 -39
rect 266 -40 267 -39
rect 267 -40 268 -39
rect 268 -40 269 -39
rect 269 -40 270 -39
rect 270 -40 271 -39
rect 271 -40 272 -39
rect 272 -40 273 -39
rect 273 -40 274 -39
rect 274 -40 275 -39
rect 275 -40 276 -39
rect 276 -40 277 -39
rect 277 -40 278 -39
rect 278 -40 279 -39
rect 279 -40 280 -39
rect 280 -40 281 -39
rect 281 -40 282 -39
rect 282 -40 283 -39
rect 283 -40 284 -39
rect 284 -40 285 -39
rect 285 -40 286 -39
rect 286 -40 287 -39
rect 287 -40 288 -39
rect 288 -40 289 -39
rect 289 -40 290 -39
rect 290 -40 291 -39
rect 291 -40 292 -39
rect 292 -40 293 -39
rect 293 -40 294 -39
rect 294 -40 295 -39
rect 295 -40 296 -39
rect 296 -40 297 -39
rect 297 -40 298 -39
rect 298 -40 299 -39
rect 299 -40 300 -39
rect 300 -40 301 -39
rect 301 -40 302 -39
rect 302 -40 303 -39
rect 303 -40 304 -39
rect 304 -40 305 -39
rect 305 -40 306 -39
rect 306 -40 307 -39
rect 307 -40 308 -39
rect 308 -40 309 -39
rect 309 -40 310 -39
rect 310 -40 311 -39
rect 311 -40 312 -39
rect 312 -40 313 -39
rect 313 -40 314 -39
rect 314 -40 315 -39
rect 315 -40 316 -39
rect 316 -40 317 -39
rect 317 -40 318 -39
rect 318 -40 319 -39
rect 319 -40 320 -39
rect 320 -40 321 -39
rect 321 -40 322 -39
rect 322 -40 323 -39
rect 323 -40 324 -39
rect 324 -40 325 -39
rect 325 -40 326 -39
rect 326 -40 327 -39
rect 327 -40 328 -39
rect 328 -40 329 -39
rect 329 -40 330 -39
rect 330 -40 331 -39
rect 331 -40 332 -39
rect 332 -40 333 -39
rect 333 -40 334 -39
rect 334 -40 335 -39
rect 335 -40 336 -39
rect 336 -40 337 -39
rect 337 -40 338 -39
rect 338 -40 339 -39
rect 339 -40 340 -39
rect 340 -40 341 -39
rect 341 -40 342 -39
rect 342 -40 343 -39
rect 343 -40 344 -39
rect 344 -40 345 -39
rect 345 -40 346 -39
rect 346 -40 347 -39
rect 347 -40 348 -39
rect 348 -40 349 -39
rect 349 -40 350 -39
rect 350 -40 351 -39
rect 351 -40 352 -39
rect 352 -40 353 -39
rect 353 -40 354 -39
rect 354 -40 355 -39
rect 355 -40 356 -39
rect 356 -40 357 -39
rect 357 -40 358 -39
rect 358 -40 359 -39
rect 359 -40 360 -39
rect 360 -40 361 -39
rect 361 -40 362 -39
rect 362 -40 363 -39
rect 363 -40 364 -39
rect 364 -40 365 -39
rect 365 -40 366 -39
rect 366 -40 367 -39
rect 367 -40 368 -39
rect 368 -40 369 -39
rect 369 -40 370 -39
rect 370 -40 371 -39
rect 371 -40 372 -39
rect 372 -40 373 -39
rect 373 -40 374 -39
rect 374 -40 375 -39
rect 375 -40 376 -39
rect 376 -40 377 -39
rect 377 -40 378 -39
rect 378 -40 379 -39
rect 379 -40 380 -39
rect 380 -40 381 -39
rect 381 -40 382 -39
rect 382 -40 383 -39
rect 383 -40 384 -39
rect 384 -40 385 -39
rect 385 -40 386 -39
rect 386 -40 387 -39
rect 387 -40 388 -39
rect 388 -40 389 -39
rect 389 -40 390 -39
rect 390 -40 391 -39
rect 391 -40 392 -39
rect 392 -40 393 -39
rect 393 -40 394 -39
rect 394 -40 395 -39
rect 395 -40 396 -39
rect 396 -40 397 -39
rect 397 -40 398 -39
rect 398 -40 399 -39
rect 399 -40 400 -39
rect 400 -40 401 -39
rect 401 -40 402 -39
rect 402 -40 403 -39
rect 403 -40 404 -39
rect 404 -40 405 -39
rect 405 -40 406 -39
rect 406 -40 407 -39
rect 407 -40 408 -39
rect 408 -40 409 -39
rect 409 -40 410 -39
rect 410 -40 411 -39
rect 411 -40 412 -39
rect 412 -40 413 -39
rect 413 -40 414 -39
rect 414 -40 415 -39
rect 415 -40 416 -39
rect 416 -40 417 -39
rect 417 -40 418 -39
rect 418 -40 419 -39
rect 419 -40 420 -39
rect 420 -40 421 -39
rect 421 -40 422 -39
rect 422 -40 423 -39
rect 423 -40 424 -39
rect 424 -40 425 -39
rect 425 -40 426 -39
rect 426 -40 427 -39
rect 427 -40 428 -39
rect 428 -40 429 -39
rect 429 -40 430 -39
rect 430 -40 431 -39
rect 431 -40 432 -39
rect 432 -40 433 -39
rect 433 -40 434 -39
rect 434 -40 435 -39
rect 435 -40 436 -39
rect 436 -40 437 -39
rect 437 -40 438 -39
rect 438 -40 439 -39
rect 439 -40 440 -39
rect 440 -40 441 -39
rect 441 -40 442 -39
rect 442 -40 443 -39
rect 443 -40 444 -39
rect 444 -40 445 -39
rect 445 -40 446 -39
rect 446 -40 447 -39
rect 447 -40 448 -39
rect 448 -40 449 -39
rect 449 -40 450 -39
rect 450 -40 451 -39
rect 451 -40 452 -39
rect 452 -40 453 -39
rect 453 -40 454 -39
rect 454 -40 455 -39
rect 455 -40 456 -39
rect 456 -40 457 -39
rect 457 -40 458 -39
rect 458 -40 459 -39
rect 459 -40 460 -39
rect 460 -40 461 -39
rect 461 -40 462 -39
rect 462 -40 463 -39
rect 463 -40 464 -39
rect 464 -40 465 -39
rect 465 -40 466 -39
rect 466 -40 467 -39
rect 467 -40 468 -39
rect 468 -40 469 -39
rect 469 -40 470 -39
rect 470 -40 471 -39
rect 471 -40 472 -39
rect 472 -40 473 -39
rect 473 -40 474 -39
rect 474 -40 475 -39
rect 475 -40 476 -39
rect 476 -40 477 -39
rect 477 -40 478 -39
rect 478 -40 479 -39
rect 479 -40 480 -39
rect 2 -41 3 -40
rect 3 -41 4 -40
rect 4 -41 5 -40
rect 5 -41 6 -40
rect 6 -41 7 -40
rect 7 -41 8 -40
rect 8 -41 9 -40
rect 9 -41 10 -40
rect 10 -41 11 -40
rect 22 -41 23 -40
rect 23 -41 24 -40
rect 24 -41 25 -40
rect 25 -41 26 -40
rect 26 -41 27 -40
rect 27 -41 28 -40
rect 28 -41 29 -40
rect 29 -41 30 -40
rect 30 -41 31 -40
rect 31 -41 32 -40
rect 32 -41 33 -40
rect 33 -41 34 -40
rect 34 -41 35 -40
rect 35 -41 36 -40
rect 36 -41 37 -40
rect 37 -41 38 -40
rect 38 -41 39 -40
rect 39 -41 40 -40
rect 40 -41 41 -40
rect 41 -41 42 -40
rect 42 -41 43 -40
rect 54 -41 55 -40
rect 55 -41 56 -40
rect 56 -41 57 -40
rect 57 -41 58 -40
rect 58 -41 59 -40
rect 59 -41 60 -40
rect 60 -41 61 -40
rect 61 -41 62 -40
rect 62 -41 63 -40
rect 63 -41 64 -40
rect 64 -41 65 -40
rect 65 -41 66 -40
rect 66 -41 67 -40
rect 67 -41 68 -40
rect 68 -41 69 -40
rect 69 -41 70 -40
rect 70 -41 71 -40
rect 71 -41 72 -40
rect 72 -41 73 -40
rect 73 -41 74 -40
rect 74 -41 75 -40
rect 86 -41 87 -40
rect 87 -41 88 -40
rect 88 -41 89 -40
rect 89 -41 90 -40
rect 90 -41 91 -40
rect 91 -41 92 -40
rect 92 -41 93 -40
rect 93 -41 94 -40
rect 94 -41 95 -40
rect 95 -41 96 -40
rect 96 -41 97 -40
rect 97 -41 98 -40
rect 98 -41 99 -40
rect 99 -41 100 -40
rect 100 -41 101 -40
rect 101 -41 102 -40
rect 102 -41 103 -40
rect 103 -41 104 -40
rect 104 -41 105 -40
rect 105 -41 106 -40
rect 106 -41 107 -40
rect 118 -41 119 -40
rect 119 -41 120 -40
rect 120 -41 121 -40
rect 121 -41 122 -40
rect 122 -41 123 -40
rect 123 -41 124 -40
rect 124 -41 125 -40
rect 125 -41 126 -40
rect 126 -41 127 -40
rect 127 -41 128 -40
rect 128 -41 129 -40
rect 129 -41 130 -40
rect 130 -41 131 -40
rect 131 -41 132 -40
rect 132 -41 133 -40
rect 133 -41 134 -40
rect 134 -41 135 -40
rect 135 -41 136 -40
rect 136 -41 137 -40
rect 137 -41 138 -40
rect 138 -41 139 -40
rect 150 -41 151 -40
rect 151 -41 152 -40
rect 152 -41 153 -40
rect 153 -41 154 -40
rect 154 -41 155 -40
rect 155 -41 156 -40
rect 156 -41 157 -40
rect 157 -41 158 -40
rect 158 -41 159 -40
rect 159 -41 160 -40
rect 160 -41 161 -40
rect 161 -41 162 -40
rect 162 -41 163 -40
rect 163 -41 164 -40
rect 164 -41 165 -40
rect 165 -41 166 -40
rect 166 -41 167 -40
rect 167 -41 168 -40
rect 168 -41 169 -40
rect 169 -41 170 -40
rect 170 -41 171 -40
rect 182 -41 183 -40
rect 183 -41 184 -40
rect 184 -41 185 -40
rect 185 -41 186 -40
rect 186 -41 187 -40
rect 187 -41 188 -40
rect 188 -41 189 -40
rect 189 -41 190 -40
rect 190 -41 191 -40
rect 191 -41 192 -40
rect 192 -41 193 -40
rect 193 -41 194 -40
rect 194 -41 195 -40
rect 195 -41 196 -40
rect 196 -41 197 -40
rect 197 -41 198 -40
rect 198 -41 199 -40
rect 199 -41 200 -40
rect 200 -41 201 -40
rect 201 -41 202 -40
rect 202 -41 203 -40
rect 203 -41 204 -40
rect 204 -41 205 -40
rect 205 -41 206 -40
rect 206 -41 207 -40
rect 207 -41 208 -40
rect 208 -41 209 -40
rect 209 -41 210 -40
rect 210 -41 211 -40
rect 211 -41 212 -40
rect 212 -41 213 -40
rect 213 -41 214 -40
rect 214 -41 215 -40
rect 215 -41 216 -40
rect 216 -41 217 -40
rect 217 -41 218 -40
rect 218 -41 219 -40
rect 219 -41 220 -40
rect 220 -41 221 -40
rect 221 -41 222 -40
rect 222 -41 223 -40
rect 223 -41 224 -40
rect 224 -41 225 -40
rect 225 -41 226 -40
rect 226 -41 227 -40
rect 227 -41 228 -40
rect 228 -41 229 -40
rect 229 -41 230 -40
rect 230 -41 231 -40
rect 231 -41 232 -40
rect 232 -41 233 -40
rect 233 -41 234 -40
rect 234 -41 235 -40
rect 235 -41 236 -40
rect 236 -41 237 -40
rect 237 -41 238 -40
rect 238 -41 239 -40
rect 239 -41 240 -40
rect 240 -41 241 -40
rect 241 -41 242 -40
rect 242 -41 243 -40
rect 243 -41 244 -40
rect 244 -41 245 -40
rect 245 -41 246 -40
rect 246 -41 247 -40
rect 247 -41 248 -40
rect 248 -41 249 -40
rect 249 -41 250 -40
rect 250 -41 251 -40
rect 251 -41 252 -40
rect 252 -41 253 -40
rect 253 -41 254 -40
rect 254 -41 255 -40
rect 255 -41 256 -40
rect 256 -41 257 -40
rect 257 -41 258 -40
rect 258 -41 259 -40
rect 259 -41 260 -40
rect 260 -41 261 -40
rect 261 -41 262 -40
rect 262 -41 263 -40
rect 263 -41 264 -40
rect 264 -41 265 -40
rect 265 -41 266 -40
rect 266 -41 267 -40
rect 267 -41 268 -40
rect 268 -41 269 -40
rect 269 -41 270 -40
rect 270 -41 271 -40
rect 271 -41 272 -40
rect 272 -41 273 -40
rect 273 -41 274 -40
rect 274 -41 275 -40
rect 275 -41 276 -40
rect 276 -41 277 -40
rect 277 -41 278 -40
rect 278 -41 279 -40
rect 279 -41 280 -40
rect 280 -41 281 -40
rect 281 -41 282 -40
rect 282 -41 283 -40
rect 283 -41 284 -40
rect 284 -41 285 -40
rect 285 -41 286 -40
rect 286 -41 287 -40
rect 287 -41 288 -40
rect 288 -41 289 -40
rect 289 -41 290 -40
rect 290 -41 291 -40
rect 291 -41 292 -40
rect 292 -41 293 -40
rect 293 -41 294 -40
rect 294 -41 295 -40
rect 295 -41 296 -40
rect 296 -41 297 -40
rect 297 -41 298 -40
rect 298 -41 299 -40
rect 299 -41 300 -40
rect 300 -41 301 -40
rect 301 -41 302 -40
rect 302 -41 303 -40
rect 303 -41 304 -40
rect 304 -41 305 -40
rect 305 -41 306 -40
rect 306 -41 307 -40
rect 307 -41 308 -40
rect 308 -41 309 -40
rect 309 -41 310 -40
rect 310 -41 311 -40
rect 311 -41 312 -40
rect 312 -41 313 -40
rect 313 -41 314 -40
rect 314 -41 315 -40
rect 315 -41 316 -40
rect 316 -41 317 -40
rect 317 -41 318 -40
rect 318 -41 319 -40
rect 319 -41 320 -40
rect 320 -41 321 -40
rect 321 -41 322 -40
rect 322 -41 323 -40
rect 323 -41 324 -40
rect 324 -41 325 -40
rect 325 -41 326 -40
rect 326 -41 327 -40
rect 327 -41 328 -40
rect 328 -41 329 -40
rect 329 -41 330 -40
rect 330 -41 331 -40
rect 331 -41 332 -40
rect 332 -41 333 -40
rect 333 -41 334 -40
rect 334 -41 335 -40
rect 335 -41 336 -40
rect 336 -41 337 -40
rect 337 -41 338 -40
rect 338 -41 339 -40
rect 339 -41 340 -40
rect 340 -41 341 -40
rect 341 -41 342 -40
rect 342 -41 343 -40
rect 343 -41 344 -40
rect 344 -41 345 -40
rect 345 -41 346 -40
rect 346 -41 347 -40
rect 347 -41 348 -40
rect 348 -41 349 -40
rect 349 -41 350 -40
rect 350 -41 351 -40
rect 351 -41 352 -40
rect 352 -41 353 -40
rect 353 -41 354 -40
rect 354 -41 355 -40
rect 355 -41 356 -40
rect 356 -41 357 -40
rect 357 -41 358 -40
rect 358 -41 359 -40
rect 359 -41 360 -40
rect 360 -41 361 -40
rect 361 -41 362 -40
rect 362 -41 363 -40
rect 363 -41 364 -40
rect 364 -41 365 -40
rect 365 -41 366 -40
rect 366 -41 367 -40
rect 367 -41 368 -40
rect 368 -41 369 -40
rect 369 -41 370 -40
rect 370 -41 371 -40
rect 371 -41 372 -40
rect 372 -41 373 -40
rect 373 -41 374 -40
rect 374 -41 375 -40
rect 375 -41 376 -40
rect 376 -41 377 -40
rect 377 -41 378 -40
rect 378 -41 379 -40
rect 379 -41 380 -40
rect 380 -41 381 -40
rect 381 -41 382 -40
rect 382 -41 383 -40
rect 383 -41 384 -40
rect 384 -41 385 -40
rect 385 -41 386 -40
rect 386 -41 387 -40
rect 387 -41 388 -40
rect 388 -41 389 -40
rect 389 -41 390 -40
rect 390 -41 391 -40
rect 391 -41 392 -40
rect 392 -41 393 -40
rect 393 -41 394 -40
rect 394 -41 395 -40
rect 395 -41 396 -40
rect 396 -41 397 -40
rect 397 -41 398 -40
rect 398 -41 399 -40
rect 399 -41 400 -40
rect 400 -41 401 -40
rect 401 -41 402 -40
rect 402 -41 403 -40
rect 403 -41 404 -40
rect 404 -41 405 -40
rect 405 -41 406 -40
rect 406 -41 407 -40
rect 407 -41 408 -40
rect 408 -41 409 -40
rect 409 -41 410 -40
rect 410 -41 411 -40
rect 411 -41 412 -40
rect 412 -41 413 -40
rect 413 -41 414 -40
rect 414 -41 415 -40
rect 415 -41 416 -40
rect 416 -41 417 -40
rect 417 -41 418 -40
rect 418 -41 419 -40
rect 419 -41 420 -40
rect 420 -41 421 -40
rect 421 -41 422 -40
rect 422 -41 423 -40
rect 423 -41 424 -40
rect 424 -41 425 -40
rect 425 -41 426 -40
rect 426 -41 427 -40
rect 427 -41 428 -40
rect 428 -41 429 -40
rect 429 -41 430 -40
rect 430 -41 431 -40
rect 431 -41 432 -40
rect 432 -41 433 -40
rect 433 -41 434 -40
rect 434 -41 435 -40
rect 435 -41 436 -40
rect 436 -41 437 -40
rect 437 -41 438 -40
rect 438 -41 439 -40
rect 439 -41 440 -40
rect 440 -41 441 -40
rect 441 -41 442 -40
rect 442 -41 443 -40
rect 443 -41 444 -40
rect 444 -41 445 -40
rect 445 -41 446 -40
rect 446 -41 447 -40
rect 447 -41 448 -40
rect 448 -41 449 -40
rect 449 -41 450 -40
rect 450 -41 451 -40
rect 451 -41 452 -40
rect 452 -41 453 -40
rect 453 -41 454 -40
rect 454 -41 455 -40
rect 455 -41 456 -40
rect 456 -41 457 -40
rect 457 -41 458 -40
rect 458 -41 459 -40
rect 459 -41 460 -40
rect 460 -41 461 -40
rect 461 -41 462 -40
rect 462 -41 463 -40
rect 463 -41 464 -40
rect 464 -41 465 -40
rect 465 -41 466 -40
rect 466 -41 467 -40
rect 467 -41 468 -40
rect 468 -41 469 -40
rect 469 -41 470 -40
rect 470 -41 471 -40
rect 471 -41 472 -40
rect 472 -41 473 -40
rect 473 -41 474 -40
rect 474 -41 475 -40
rect 475 -41 476 -40
rect 476 -41 477 -40
rect 477 -41 478 -40
rect 478 -41 479 -40
rect 479 -41 480 -40
rect 2 -42 3 -41
rect 3 -42 4 -41
rect 4 -42 5 -41
rect 5 -42 6 -41
rect 6 -42 7 -41
rect 7 -42 8 -41
rect 8 -42 9 -41
rect 9 -42 10 -41
rect 10 -42 11 -41
rect 11 -42 12 -41
rect 21 -42 22 -41
rect 22 -42 23 -41
rect 23 -42 24 -41
rect 24 -42 25 -41
rect 25 -42 26 -41
rect 26 -42 27 -41
rect 27 -42 28 -41
rect 28 -42 29 -41
rect 29 -42 30 -41
rect 30 -42 31 -41
rect 31 -42 32 -41
rect 32 -42 33 -41
rect 33 -42 34 -41
rect 34 -42 35 -41
rect 35 -42 36 -41
rect 36 -42 37 -41
rect 37 -42 38 -41
rect 38 -42 39 -41
rect 39 -42 40 -41
rect 40 -42 41 -41
rect 41 -42 42 -41
rect 42 -42 43 -41
rect 43 -42 44 -41
rect 53 -42 54 -41
rect 54 -42 55 -41
rect 55 -42 56 -41
rect 56 -42 57 -41
rect 57 -42 58 -41
rect 58 -42 59 -41
rect 59 -42 60 -41
rect 60 -42 61 -41
rect 61 -42 62 -41
rect 62 -42 63 -41
rect 63 -42 64 -41
rect 64 -42 65 -41
rect 65 -42 66 -41
rect 66 -42 67 -41
rect 67 -42 68 -41
rect 68 -42 69 -41
rect 69 -42 70 -41
rect 70 -42 71 -41
rect 71 -42 72 -41
rect 72 -42 73 -41
rect 73 -42 74 -41
rect 74 -42 75 -41
rect 75 -42 76 -41
rect 85 -42 86 -41
rect 86 -42 87 -41
rect 87 -42 88 -41
rect 88 -42 89 -41
rect 89 -42 90 -41
rect 90 -42 91 -41
rect 91 -42 92 -41
rect 92 -42 93 -41
rect 93 -42 94 -41
rect 94 -42 95 -41
rect 95 -42 96 -41
rect 96 -42 97 -41
rect 97 -42 98 -41
rect 98 -42 99 -41
rect 99 -42 100 -41
rect 100 -42 101 -41
rect 101 -42 102 -41
rect 102 -42 103 -41
rect 103 -42 104 -41
rect 104 -42 105 -41
rect 105 -42 106 -41
rect 106 -42 107 -41
rect 107 -42 108 -41
rect 117 -42 118 -41
rect 118 -42 119 -41
rect 119 -42 120 -41
rect 120 -42 121 -41
rect 121 -42 122 -41
rect 122 -42 123 -41
rect 123 -42 124 -41
rect 124 -42 125 -41
rect 125 -42 126 -41
rect 126 -42 127 -41
rect 127 -42 128 -41
rect 128 -42 129 -41
rect 129 -42 130 -41
rect 130 -42 131 -41
rect 131 -42 132 -41
rect 132 -42 133 -41
rect 133 -42 134 -41
rect 134 -42 135 -41
rect 135 -42 136 -41
rect 136 -42 137 -41
rect 137 -42 138 -41
rect 138 -42 139 -41
rect 139 -42 140 -41
rect 149 -42 150 -41
rect 150 -42 151 -41
rect 151 -42 152 -41
rect 152 -42 153 -41
rect 153 -42 154 -41
rect 154 -42 155 -41
rect 155 -42 156 -41
rect 156 -42 157 -41
rect 157 -42 158 -41
rect 158 -42 159 -41
rect 159 -42 160 -41
rect 160 -42 161 -41
rect 161 -42 162 -41
rect 162 -42 163 -41
rect 163 -42 164 -41
rect 164 -42 165 -41
rect 165 -42 166 -41
rect 166 -42 167 -41
rect 167 -42 168 -41
rect 168 -42 169 -41
rect 169 -42 170 -41
rect 170 -42 171 -41
rect 171 -42 172 -41
rect 181 -42 182 -41
rect 182 -42 183 -41
rect 183 -42 184 -41
rect 184 -42 185 -41
rect 185 -42 186 -41
rect 186 -42 187 -41
rect 187 -42 188 -41
rect 188 -42 189 -41
rect 189 -42 190 -41
rect 190 -42 191 -41
rect 191 -42 192 -41
rect 192 -42 193 -41
rect 193 -42 194 -41
rect 194 -42 195 -41
rect 195 -42 196 -41
rect 196 -42 197 -41
rect 197 -42 198 -41
rect 198 -42 199 -41
rect 199 -42 200 -41
rect 200 -42 201 -41
rect 201 -42 202 -41
rect 202 -42 203 -41
rect 203 -42 204 -41
rect 204 -42 205 -41
rect 205 -42 206 -41
rect 206 -42 207 -41
rect 207 -42 208 -41
rect 208 -42 209 -41
rect 209 -42 210 -41
rect 210 -42 211 -41
rect 211 -42 212 -41
rect 212 -42 213 -41
rect 213 -42 214 -41
rect 214 -42 215 -41
rect 215 -42 216 -41
rect 216 -42 217 -41
rect 217 -42 218 -41
rect 218 -42 219 -41
rect 219 -42 220 -41
rect 220 -42 221 -41
rect 221 -42 222 -41
rect 222 -42 223 -41
rect 223 -42 224 -41
rect 224 -42 225 -41
rect 225 -42 226 -41
rect 226 -42 227 -41
rect 227 -42 228 -41
rect 228 -42 229 -41
rect 229 -42 230 -41
rect 230 -42 231 -41
rect 231 -42 232 -41
rect 232 -42 233 -41
rect 233 -42 234 -41
rect 234 -42 235 -41
rect 235 -42 236 -41
rect 236 -42 237 -41
rect 237 -42 238 -41
rect 238 -42 239 -41
rect 239 -42 240 -41
rect 240 -42 241 -41
rect 241 -42 242 -41
rect 242 -42 243 -41
rect 243 -42 244 -41
rect 244 -42 245 -41
rect 245 -42 246 -41
rect 246 -42 247 -41
rect 247 -42 248 -41
rect 248 -42 249 -41
rect 249 -42 250 -41
rect 250 -42 251 -41
rect 251 -42 252 -41
rect 252 -42 253 -41
rect 253 -42 254 -41
rect 254 -42 255 -41
rect 255 -42 256 -41
rect 256 -42 257 -41
rect 257 -42 258 -41
rect 258 -42 259 -41
rect 259 -42 260 -41
rect 260 -42 261 -41
rect 261 -42 262 -41
rect 262 -42 263 -41
rect 263 -42 264 -41
rect 264 -42 265 -41
rect 265 -42 266 -41
rect 266 -42 267 -41
rect 267 -42 268 -41
rect 268 -42 269 -41
rect 269 -42 270 -41
rect 270 -42 271 -41
rect 271 -42 272 -41
rect 272 -42 273 -41
rect 273 -42 274 -41
rect 274 -42 275 -41
rect 275 -42 276 -41
rect 276 -42 277 -41
rect 277 -42 278 -41
rect 278 -42 279 -41
rect 279 -42 280 -41
rect 280 -42 281 -41
rect 281 -42 282 -41
rect 282 -42 283 -41
rect 283 -42 284 -41
rect 284 -42 285 -41
rect 285 -42 286 -41
rect 286 -42 287 -41
rect 287 -42 288 -41
rect 288 -42 289 -41
rect 289 -42 290 -41
rect 290 -42 291 -41
rect 291 -42 292 -41
rect 292 -42 293 -41
rect 293 -42 294 -41
rect 294 -42 295 -41
rect 295 -42 296 -41
rect 296 -42 297 -41
rect 297 -42 298 -41
rect 298 -42 299 -41
rect 299 -42 300 -41
rect 300 -42 301 -41
rect 301 -42 302 -41
rect 302 -42 303 -41
rect 303 -42 304 -41
rect 304 -42 305 -41
rect 305 -42 306 -41
rect 306 -42 307 -41
rect 307 -42 308 -41
rect 308 -42 309 -41
rect 309 -42 310 -41
rect 310 -42 311 -41
rect 311 -42 312 -41
rect 312 -42 313 -41
rect 313 -42 314 -41
rect 314 -42 315 -41
rect 315 -42 316 -41
rect 316 -42 317 -41
rect 317 -42 318 -41
rect 318 -42 319 -41
rect 319 -42 320 -41
rect 320 -42 321 -41
rect 321 -42 322 -41
rect 322 -42 323 -41
rect 323 -42 324 -41
rect 324 -42 325 -41
rect 325 -42 326 -41
rect 326 -42 327 -41
rect 327 -42 328 -41
rect 328 -42 329 -41
rect 329 -42 330 -41
rect 330 -42 331 -41
rect 331 -42 332 -41
rect 332 -42 333 -41
rect 333 -42 334 -41
rect 334 -42 335 -41
rect 335 -42 336 -41
rect 336 -42 337 -41
rect 337 -42 338 -41
rect 338 -42 339 -41
rect 339 -42 340 -41
rect 340 -42 341 -41
rect 341 -42 342 -41
rect 342 -42 343 -41
rect 343 -42 344 -41
rect 344 -42 345 -41
rect 345 -42 346 -41
rect 346 -42 347 -41
rect 347 -42 348 -41
rect 348 -42 349 -41
rect 349 -42 350 -41
rect 350 -42 351 -41
rect 351 -42 352 -41
rect 352 -42 353 -41
rect 353 -42 354 -41
rect 354 -42 355 -41
rect 355 -42 356 -41
rect 356 -42 357 -41
rect 357 -42 358 -41
rect 358 -42 359 -41
rect 359 -42 360 -41
rect 360 -42 361 -41
rect 361 -42 362 -41
rect 362 -42 363 -41
rect 363 -42 364 -41
rect 364 -42 365 -41
rect 365 -42 366 -41
rect 366 -42 367 -41
rect 367 -42 368 -41
rect 368 -42 369 -41
rect 369 -42 370 -41
rect 370 -42 371 -41
rect 371 -42 372 -41
rect 372 -42 373 -41
rect 373 -42 374 -41
rect 374 -42 375 -41
rect 375 -42 376 -41
rect 376 -42 377 -41
rect 377 -42 378 -41
rect 378 -42 379 -41
rect 379 -42 380 -41
rect 380 -42 381 -41
rect 381 -42 382 -41
rect 382 -42 383 -41
rect 383 -42 384 -41
rect 384 -42 385 -41
rect 385 -42 386 -41
rect 386 -42 387 -41
rect 387 -42 388 -41
rect 388 -42 389 -41
rect 389 -42 390 -41
rect 390 -42 391 -41
rect 391 -42 392 -41
rect 392 -42 393 -41
rect 393 -42 394 -41
rect 394 -42 395 -41
rect 395 -42 396 -41
rect 396 -42 397 -41
rect 397 -42 398 -41
rect 398 -42 399 -41
rect 399 -42 400 -41
rect 400 -42 401 -41
rect 401 -42 402 -41
rect 402 -42 403 -41
rect 403 -42 404 -41
rect 404 -42 405 -41
rect 405 -42 406 -41
rect 406 -42 407 -41
rect 407 -42 408 -41
rect 408 -42 409 -41
rect 409 -42 410 -41
rect 410 -42 411 -41
rect 411 -42 412 -41
rect 412 -42 413 -41
rect 413 -42 414 -41
rect 414 -42 415 -41
rect 415 -42 416 -41
rect 416 -42 417 -41
rect 417 -42 418 -41
rect 418 -42 419 -41
rect 419 -42 420 -41
rect 420 -42 421 -41
rect 421 -42 422 -41
rect 422 -42 423 -41
rect 423 -42 424 -41
rect 424 -42 425 -41
rect 425 -42 426 -41
rect 426 -42 427 -41
rect 427 -42 428 -41
rect 428 -42 429 -41
rect 429 -42 430 -41
rect 430 -42 431 -41
rect 431 -42 432 -41
rect 432 -42 433 -41
rect 433 -42 434 -41
rect 434 -42 435 -41
rect 435 -42 436 -41
rect 436 -42 437 -41
rect 437 -42 438 -41
rect 438 -42 439 -41
rect 439 -42 440 -41
rect 440 -42 441 -41
rect 441 -42 442 -41
rect 442 -42 443 -41
rect 443 -42 444 -41
rect 444 -42 445 -41
rect 445 -42 446 -41
rect 446 -42 447 -41
rect 447 -42 448 -41
rect 448 -42 449 -41
rect 449 -42 450 -41
rect 450 -42 451 -41
rect 451 -42 452 -41
rect 452 -42 453 -41
rect 453 -42 454 -41
rect 454 -42 455 -41
rect 455 -42 456 -41
rect 456 -42 457 -41
rect 457 -42 458 -41
rect 458 -42 459 -41
rect 459 -42 460 -41
rect 460 -42 461 -41
rect 461 -42 462 -41
rect 462 -42 463 -41
rect 463 -42 464 -41
rect 464 -42 465 -41
rect 465 -42 466 -41
rect 466 -42 467 -41
rect 467 -42 468 -41
rect 468 -42 469 -41
rect 469 -42 470 -41
rect 470 -42 471 -41
rect 471 -42 472 -41
rect 472 -42 473 -41
rect 473 -42 474 -41
rect 474 -42 475 -41
rect 475 -42 476 -41
rect 476 -42 477 -41
rect 477 -42 478 -41
rect 478 -42 479 -41
rect 479 -42 480 -41
rect 2 -43 3 -42
rect 3 -43 4 -42
rect 4 -43 5 -42
rect 5 -43 6 -42
rect 6 -43 7 -42
rect 7 -43 8 -42
rect 8 -43 9 -42
rect 9 -43 10 -42
rect 10 -43 11 -42
rect 11 -43 12 -42
rect 21 -43 22 -42
rect 22 -43 23 -42
rect 23 -43 24 -42
rect 24 -43 25 -42
rect 25 -43 26 -42
rect 26 -43 27 -42
rect 27 -43 28 -42
rect 28 -43 29 -42
rect 29 -43 30 -42
rect 30 -43 31 -42
rect 31 -43 32 -42
rect 32 -43 33 -42
rect 33 -43 34 -42
rect 34 -43 35 -42
rect 35 -43 36 -42
rect 36 -43 37 -42
rect 37 -43 38 -42
rect 38 -43 39 -42
rect 39 -43 40 -42
rect 40 -43 41 -42
rect 41 -43 42 -42
rect 42 -43 43 -42
rect 43 -43 44 -42
rect 53 -43 54 -42
rect 54 -43 55 -42
rect 55 -43 56 -42
rect 56 -43 57 -42
rect 57 -43 58 -42
rect 58 -43 59 -42
rect 59 -43 60 -42
rect 60 -43 61 -42
rect 61 -43 62 -42
rect 62 -43 63 -42
rect 63 -43 64 -42
rect 64 -43 65 -42
rect 65 -43 66 -42
rect 66 -43 67 -42
rect 67 -43 68 -42
rect 68 -43 69 -42
rect 69 -43 70 -42
rect 70 -43 71 -42
rect 71 -43 72 -42
rect 72 -43 73 -42
rect 73 -43 74 -42
rect 74 -43 75 -42
rect 75 -43 76 -42
rect 85 -43 86 -42
rect 86 -43 87 -42
rect 87 -43 88 -42
rect 88 -43 89 -42
rect 89 -43 90 -42
rect 90 -43 91 -42
rect 91 -43 92 -42
rect 92 -43 93 -42
rect 93 -43 94 -42
rect 94 -43 95 -42
rect 95 -43 96 -42
rect 96 -43 97 -42
rect 97 -43 98 -42
rect 98 -43 99 -42
rect 99 -43 100 -42
rect 100 -43 101 -42
rect 101 -43 102 -42
rect 102 -43 103 -42
rect 103 -43 104 -42
rect 104 -43 105 -42
rect 105 -43 106 -42
rect 106 -43 107 -42
rect 107 -43 108 -42
rect 117 -43 118 -42
rect 118 -43 119 -42
rect 119 -43 120 -42
rect 120 -43 121 -42
rect 121 -43 122 -42
rect 122 -43 123 -42
rect 123 -43 124 -42
rect 124 -43 125 -42
rect 125 -43 126 -42
rect 126 -43 127 -42
rect 127 -43 128 -42
rect 128 -43 129 -42
rect 129 -43 130 -42
rect 130 -43 131 -42
rect 131 -43 132 -42
rect 132 -43 133 -42
rect 133 -43 134 -42
rect 134 -43 135 -42
rect 135 -43 136 -42
rect 136 -43 137 -42
rect 137 -43 138 -42
rect 138 -43 139 -42
rect 139 -43 140 -42
rect 149 -43 150 -42
rect 150 -43 151 -42
rect 151 -43 152 -42
rect 152 -43 153 -42
rect 153 -43 154 -42
rect 154 -43 155 -42
rect 155 -43 156 -42
rect 156 -43 157 -42
rect 157 -43 158 -42
rect 158 -43 159 -42
rect 159 -43 160 -42
rect 160 -43 161 -42
rect 161 -43 162 -42
rect 162 -43 163 -42
rect 163 -43 164 -42
rect 164 -43 165 -42
rect 165 -43 166 -42
rect 166 -43 167 -42
rect 167 -43 168 -42
rect 168 -43 169 -42
rect 169 -43 170 -42
rect 170 -43 171 -42
rect 171 -43 172 -42
rect 181 -43 182 -42
rect 182 -43 183 -42
rect 183 -43 184 -42
rect 184 -43 185 -42
rect 185 -43 186 -42
rect 186 -43 187 -42
rect 187 -43 188 -42
rect 188 -43 189 -42
rect 189 -43 190 -42
rect 190 -43 191 -42
rect 191 -43 192 -42
rect 192 -43 193 -42
rect 193 -43 194 -42
rect 194 -43 195 -42
rect 195 -43 196 -42
rect 196 -43 197 -42
rect 197 -43 198 -42
rect 198 -43 199 -42
rect 199 -43 200 -42
rect 200 -43 201 -42
rect 201 -43 202 -42
rect 202 -43 203 -42
rect 203 -43 204 -42
rect 204 -43 205 -42
rect 205 -43 206 -42
rect 206 -43 207 -42
rect 207 -43 208 -42
rect 208 -43 209 -42
rect 209 -43 210 -42
rect 210 -43 211 -42
rect 211 -43 212 -42
rect 212 -43 213 -42
rect 213 -43 214 -42
rect 214 -43 215 -42
rect 215 -43 216 -42
rect 216 -43 217 -42
rect 217 -43 218 -42
rect 218 -43 219 -42
rect 219 -43 220 -42
rect 220 -43 221 -42
rect 221 -43 222 -42
rect 222 -43 223 -42
rect 223 -43 224 -42
rect 224 -43 225 -42
rect 225 -43 226 -42
rect 226 -43 227 -42
rect 227 -43 228 -42
rect 228 -43 229 -42
rect 229 -43 230 -42
rect 230 -43 231 -42
rect 231 -43 232 -42
rect 232 -43 233 -42
rect 233 -43 234 -42
rect 234 -43 235 -42
rect 235 -43 236 -42
rect 236 -43 237 -42
rect 237 -43 238 -42
rect 238 -43 239 -42
rect 239 -43 240 -42
rect 240 -43 241 -42
rect 241 -43 242 -42
rect 242 -43 243 -42
rect 243 -43 244 -42
rect 244 -43 245 -42
rect 245 -43 246 -42
rect 246 -43 247 -42
rect 247 -43 248 -42
rect 248 -43 249 -42
rect 249 -43 250 -42
rect 250 -43 251 -42
rect 251 -43 252 -42
rect 252 -43 253 -42
rect 253 -43 254 -42
rect 254 -43 255 -42
rect 255 -43 256 -42
rect 256 -43 257 -42
rect 257 -43 258 -42
rect 258 -43 259 -42
rect 259 -43 260 -42
rect 260 -43 261 -42
rect 261 -43 262 -42
rect 262 -43 263 -42
rect 263 -43 264 -42
rect 264 -43 265 -42
rect 265 -43 266 -42
rect 266 -43 267 -42
rect 267 -43 268 -42
rect 268 -43 269 -42
rect 269 -43 270 -42
rect 270 -43 271 -42
rect 271 -43 272 -42
rect 272 -43 273 -42
rect 273 -43 274 -42
rect 274 -43 275 -42
rect 275 -43 276 -42
rect 276 -43 277 -42
rect 277 -43 278 -42
rect 278 -43 279 -42
rect 279 -43 280 -42
rect 280 -43 281 -42
rect 281 -43 282 -42
rect 282 -43 283 -42
rect 283 -43 284 -42
rect 284 -43 285 -42
rect 285 -43 286 -42
rect 286 -43 287 -42
rect 287 -43 288 -42
rect 288 -43 289 -42
rect 289 -43 290 -42
rect 290 -43 291 -42
rect 291 -43 292 -42
rect 292 -43 293 -42
rect 293 -43 294 -42
rect 294 -43 295 -42
rect 295 -43 296 -42
rect 296 -43 297 -42
rect 297 -43 298 -42
rect 298 -43 299 -42
rect 299 -43 300 -42
rect 300 -43 301 -42
rect 301 -43 302 -42
rect 302 -43 303 -42
rect 303 -43 304 -42
rect 304 -43 305 -42
rect 305 -43 306 -42
rect 306 -43 307 -42
rect 307 -43 308 -42
rect 308 -43 309 -42
rect 309 -43 310 -42
rect 310 -43 311 -42
rect 311 -43 312 -42
rect 312 -43 313 -42
rect 313 -43 314 -42
rect 314 -43 315 -42
rect 315 -43 316 -42
rect 316 -43 317 -42
rect 317 -43 318 -42
rect 318 -43 319 -42
rect 319 -43 320 -42
rect 320 -43 321 -42
rect 321 -43 322 -42
rect 322 -43 323 -42
rect 323 -43 324 -42
rect 324 -43 325 -42
rect 325 -43 326 -42
rect 326 -43 327 -42
rect 327 -43 328 -42
rect 328 -43 329 -42
rect 329 -43 330 -42
rect 330 -43 331 -42
rect 331 -43 332 -42
rect 332 -43 333 -42
rect 333 -43 334 -42
rect 334 -43 335 -42
rect 335 -43 336 -42
rect 336 -43 337 -42
rect 337 -43 338 -42
rect 338 -43 339 -42
rect 339 -43 340 -42
rect 340 -43 341 -42
rect 341 -43 342 -42
rect 342 -43 343 -42
rect 343 -43 344 -42
rect 344 -43 345 -42
rect 345 -43 346 -42
rect 346 -43 347 -42
rect 347 -43 348 -42
rect 348 -43 349 -42
rect 349 -43 350 -42
rect 350 -43 351 -42
rect 351 -43 352 -42
rect 352 -43 353 -42
rect 353 -43 354 -42
rect 354 -43 355 -42
rect 355 -43 356 -42
rect 356 -43 357 -42
rect 357 -43 358 -42
rect 358 -43 359 -42
rect 359 -43 360 -42
rect 360 -43 361 -42
rect 361 -43 362 -42
rect 362 -43 363 -42
rect 363 -43 364 -42
rect 364 -43 365 -42
rect 365 -43 366 -42
rect 366 -43 367 -42
rect 367 -43 368 -42
rect 368 -43 369 -42
rect 369 -43 370 -42
rect 370 -43 371 -42
rect 371 -43 372 -42
rect 372 -43 373 -42
rect 373 -43 374 -42
rect 374 -43 375 -42
rect 375 -43 376 -42
rect 376 -43 377 -42
rect 377 -43 378 -42
rect 378 -43 379 -42
rect 379 -43 380 -42
rect 380 -43 381 -42
rect 381 -43 382 -42
rect 382 -43 383 -42
rect 383 -43 384 -42
rect 384 -43 385 -42
rect 385 -43 386 -42
rect 386 -43 387 -42
rect 387 -43 388 -42
rect 388 -43 389 -42
rect 389 -43 390 -42
rect 390 -43 391 -42
rect 391 -43 392 -42
rect 392 -43 393 -42
rect 393 -43 394 -42
rect 394 -43 395 -42
rect 395 -43 396 -42
rect 396 -43 397 -42
rect 397 -43 398 -42
rect 398 -43 399 -42
rect 399 -43 400 -42
rect 400 -43 401 -42
rect 401 -43 402 -42
rect 402 -43 403 -42
rect 403 -43 404 -42
rect 404 -43 405 -42
rect 405 -43 406 -42
rect 406 -43 407 -42
rect 407 -43 408 -42
rect 408 -43 409 -42
rect 409 -43 410 -42
rect 410 -43 411 -42
rect 411 -43 412 -42
rect 412 -43 413 -42
rect 413 -43 414 -42
rect 414 -43 415 -42
rect 415 -43 416 -42
rect 416 -43 417 -42
rect 417 -43 418 -42
rect 418 -43 419 -42
rect 419 -43 420 -42
rect 420 -43 421 -42
rect 421 -43 422 -42
rect 422 -43 423 -42
rect 423 -43 424 -42
rect 424 -43 425 -42
rect 425 -43 426 -42
rect 426 -43 427 -42
rect 427 -43 428 -42
rect 428 -43 429 -42
rect 429 -43 430 -42
rect 430 -43 431 -42
rect 431 -43 432 -42
rect 432 -43 433 -42
rect 433 -43 434 -42
rect 434 -43 435 -42
rect 435 -43 436 -42
rect 436 -43 437 -42
rect 437 -43 438 -42
rect 438 -43 439 -42
rect 439 -43 440 -42
rect 440 -43 441 -42
rect 441 -43 442 -42
rect 442 -43 443 -42
rect 443 -43 444 -42
rect 444 -43 445 -42
rect 445 -43 446 -42
rect 446 -43 447 -42
rect 447 -43 448 -42
rect 448 -43 449 -42
rect 449 -43 450 -42
rect 450 -43 451 -42
rect 451 -43 452 -42
rect 452 -43 453 -42
rect 453 -43 454 -42
rect 454 -43 455 -42
rect 455 -43 456 -42
rect 456 -43 457 -42
rect 457 -43 458 -42
rect 458 -43 459 -42
rect 459 -43 460 -42
rect 460 -43 461 -42
rect 461 -43 462 -42
rect 462 -43 463 -42
rect 463 -43 464 -42
rect 464 -43 465 -42
rect 465 -43 466 -42
rect 466 -43 467 -42
rect 467 -43 468 -42
rect 468 -43 469 -42
rect 469 -43 470 -42
rect 470 -43 471 -42
rect 471 -43 472 -42
rect 472 -43 473 -42
rect 473 -43 474 -42
rect 474 -43 475 -42
rect 475 -43 476 -42
rect 476 -43 477 -42
rect 477 -43 478 -42
rect 478 -43 479 -42
rect 479 -43 480 -42
rect 2 -44 3 -43
rect 3 -44 4 -43
rect 4 -44 5 -43
rect 5 -44 6 -43
rect 6 -44 7 -43
rect 7 -44 8 -43
rect 8 -44 9 -43
rect 9 -44 10 -43
rect 10 -44 11 -43
rect 11 -44 12 -43
rect 21 -44 22 -43
rect 22 -44 23 -43
rect 23 -44 24 -43
rect 24 -44 25 -43
rect 25 -44 26 -43
rect 26 -44 27 -43
rect 27 -44 28 -43
rect 28 -44 29 -43
rect 29 -44 30 -43
rect 30 -44 31 -43
rect 31 -44 32 -43
rect 32 -44 33 -43
rect 33 -44 34 -43
rect 34 -44 35 -43
rect 35 -44 36 -43
rect 36 -44 37 -43
rect 37 -44 38 -43
rect 38 -44 39 -43
rect 39 -44 40 -43
rect 40 -44 41 -43
rect 41 -44 42 -43
rect 42 -44 43 -43
rect 43 -44 44 -43
rect 53 -44 54 -43
rect 54 -44 55 -43
rect 55 -44 56 -43
rect 56 -44 57 -43
rect 57 -44 58 -43
rect 58 -44 59 -43
rect 59 -44 60 -43
rect 60 -44 61 -43
rect 61 -44 62 -43
rect 62 -44 63 -43
rect 63 -44 64 -43
rect 64 -44 65 -43
rect 65 -44 66 -43
rect 66 -44 67 -43
rect 67 -44 68 -43
rect 68 -44 69 -43
rect 69 -44 70 -43
rect 70 -44 71 -43
rect 71 -44 72 -43
rect 72 -44 73 -43
rect 73 -44 74 -43
rect 74 -44 75 -43
rect 75 -44 76 -43
rect 85 -44 86 -43
rect 86 -44 87 -43
rect 87 -44 88 -43
rect 88 -44 89 -43
rect 89 -44 90 -43
rect 90 -44 91 -43
rect 91 -44 92 -43
rect 92 -44 93 -43
rect 93 -44 94 -43
rect 94 -44 95 -43
rect 95 -44 96 -43
rect 96 -44 97 -43
rect 97 -44 98 -43
rect 98 -44 99 -43
rect 99 -44 100 -43
rect 100 -44 101 -43
rect 101 -44 102 -43
rect 102 -44 103 -43
rect 103 -44 104 -43
rect 104 -44 105 -43
rect 105 -44 106 -43
rect 106 -44 107 -43
rect 107 -44 108 -43
rect 117 -44 118 -43
rect 118 -44 119 -43
rect 119 -44 120 -43
rect 120 -44 121 -43
rect 121 -44 122 -43
rect 122 -44 123 -43
rect 123 -44 124 -43
rect 124 -44 125 -43
rect 125 -44 126 -43
rect 126 -44 127 -43
rect 127 -44 128 -43
rect 128 -44 129 -43
rect 129 -44 130 -43
rect 130 -44 131 -43
rect 131 -44 132 -43
rect 132 -44 133 -43
rect 133 -44 134 -43
rect 134 -44 135 -43
rect 135 -44 136 -43
rect 136 -44 137 -43
rect 137 -44 138 -43
rect 138 -44 139 -43
rect 139 -44 140 -43
rect 149 -44 150 -43
rect 150 -44 151 -43
rect 151 -44 152 -43
rect 152 -44 153 -43
rect 153 -44 154 -43
rect 154 -44 155 -43
rect 155 -44 156 -43
rect 156 -44 157 -43
rect 157 -44 158 -43
rect 158 -44 159 -43
rect 159 -44 160 -43
rect 160 -44 161 -43
rect 161 -44 162 -43
rect 162 -44 163 -43
rect 163 -44 164 -43
rect 164 -44 165 -43
rect 165 -44 166 -43
rect 166 -44 167 -43
rect 167 -44 168 -43
rect 168 -44 169 -43
rect 169 -44 170 -43
rect 170 -44 171 -43
rect 171 -44 172 -43
rect 181 -44 182 -43
rect 182 -44 183 -43
rect 183 -44 184 -43
rect 184 -44 185 -43
rect 185 -44 186 -43
rect 186 -44 187 -43
rect 187 -44 188 -43
rect 188 -44 189 -43
rect 189 -44 190 -43
rect 190 -44 191 -43
rect 191 -44 192 -43
rect 192 -44 193 -43
rect 193 -44 194 -43
rect 194 -44 195 -43
rect 195 -44 196 -43
rect 196 -44 197 -43
rect 197 -44 198 -43
rect 198 -44 199 -43
rect 199 -44 200 -43
rect 200 -44 201 -43
rect 201 -44 202 -43
rect 202 -44 203 -43
rect 203 -44 204 -43
rect 204 -44 205 -43
rect 205 -44 206 -43
rect 206 -44 207 -43
rect 207 -44 208 -43
rect 208 -44 209 -43
rect 209 -44 210 -43
rect 210 -44 211 -43
rect 211 -44 212 -43
rect 212 -44 213 -43
rect 213 -44 214 -43
rect 214 -44 215 -43
rect 215 -44 216 -43
rect 216 -44 217 -43
rect 217 -44 218 -43
rect 218 -44 219 -43
rect 219 -44 220 -43
rect 220 -44 221 -43
rect 221 -44 222 -43
rect 222 -44 223 -43
rect 223 -44 224 -43
rect 224 -44 225 -43
rect 225 -44 226 -43
rect 226 -44 227 -43
rect 227 -44 228 -43
rect 228 -44 229 -43
rect 229 -44 230 -43
rect 230 -44 231 -43
rect 231 -44 232 -43
rect 232 -44 233 -43
rect 233 -44 234 -43
rect 234 -44 235 -43
rect 235 -44 236 -43
rect 236 -44 237 -43
rect 237 -44 238 -43
rect 238 -44 239 -43
rect 239 -44 240 -43
rect 240 -44 241 -43
rect 241 -44 242 -43
rect 242 -44 243 -43
rect 243 -44 244 -43
rect 244 -44 245 -43
rect 245 -44 246 -43
rect 246 -44 247 -43
rect 247 -44 248 -43
rect 248 -44 249 -43
rect 249 -44 250 -43
rect 250 -44 251 -43
rect 251 -44 252 -43
rect 252 -44 253 -43
rect 253 -44 254 -43
rect 254 -44 255 -43
rect 255 -44 256 -43
rect 256 -44 257 -43
rect 257 -44 258 -43
rect 258 -44 259 -43
rect 259 -44 260 -43
rect 260 -44 261 -43
rect 261 -44 262 -43
rect 262 -44 263 -43
rect 263 -44 264 -43
rect 264 -44 265 -43
rect 265 -44 266 -43
rect 266 -44 267 -43
rect 267 -44 268 -43
rect 268 -44 269 -43
rect 269 -44 270 -43
rect 270 -44 271 -43
rect 271 -44 272 -43
rect 272 -44 273 -43
rect 273 -44 274 -43
rect 274 -44 275 -43
rect 275 -44 276 -43
rect 276 -44 277 -43
rect 277 -44 278 -43
rect 278 -44 279 -43
rect 279 -44 280 -43
rect 280 -44 281 -43
rect 281 -44 282 -43
rect 282 -44 283 -43
rect 283 -44 284 -43
rect 284 -44 285 -43
rect 285 -44 286 -43
rect 286 -44 287 -43
rect 287 -44 288 -43
rect 288 -44 289 -43
rect 289 -44 290 -43
rect 290 -44 291 -43
rect 291 -44 292 -43
rect 292 -44 293 -43
rect 293 -44 294 -43
rect 294 -44 295 -43
rect 295 -44 296 -43
rect 296 -44 297 -43
rect 297 -44 298 -43
rect 298 -44 299 -43
rect 299 -44 300 -43
rect 300 -44 301 -43
rect 301 -44 302 -43
rect 302 -44 303 -43
rect 303 -44 304 -43
rect 304 -44 305 -43
rect 305 -44 306 -43
rect 306 -44 307 -43
rect 307 -44 308 -43
rect 308 -44 309 -43
rect 309 -44 310 -43
rect 310 -44 311 -43
rect 311 -44 312 -43
rect 312 -44 313 -43
rect 313 -44 314 -43
rect 314 -44 315 -43
rect 315 -44 316 -43
rect 316 -44 317 -43
rect 317 -44 318 -43
rect 318 -44 319 -43
rect 319 -44 320 -43
rect 320 -44 321 -43
rect 321 -44 322 -43
rect 322 -44 323 -43
rect 323 -44 324 -43
rect 324 -44 325 -43
rect 325 -44 326 -43
rect 326 -44 327 -43
rect 327 -44 328 -43
rect 328 -44 329 -43
rect 329 -44 330 -43
rect 330 -44 331 -43
rect 331 -44 332 -43
rect 332 -44 333 -43
rect 333 -44 334 -43
rect 334 -44 335 -43
rect 335 -44 336 -43
rect 336 -44 337 -43
rect 337 -44 338 -43
rect 338 -44 339 -43
rect 339 -44 340 -43
rect 340 -44 341 -43
rect 341 -44 342 -43
rect 342 -44 343 -43
rect 343 -44 344 -43
rect 344 -44 345 -43
rect 345 -44 346 -43
rect 346 -44 347 -43
rect 347 -44 348 -43
rect 348 -44 349 -43
rect 349 -44 350 -43
rect 350 -44 351 -43
rect 351 -44 352 -43
rect 352 -44 353 -43
rect 353 -44 354 -43
rect 354 -44 355 -43
rect 355 -44 356 -43
rect 356 -44 357 -43
rect 357 -44 358 -43
rect 358 -44 359 -43
rect 359 -44 360 -43
rect 360 -44 361 -43
rect 361 -44 362 -43
rect 362 -44 363 -43
rect 363 -44 364 -43
rect 364 -44 365 -43
rect 365 -44 366 -43
rect 366 -44 367 -43
rect 367 -44 368 -43
rect 368 -44 369 -43
rect 369 -44 370 -43
rect 370 -44 371 -43
rect 371 -44 372 -43
rect 372 -44 373 -43
rect 373 -44 374 -43
rect 374 -44 375 -43
rect 375 -44 376 -43
rect 376 -44 377 -43
rect 377 -44 378 -43
rect 378 -44 379 -43
rect 379 -44 380 -43
rect 380 -44 381 -43
rect 381 -44 382 -43
rect 382 -44 383 -43
rect 383 -44 384 -43
rect 384 -44 385 -43
rect 385 -44 386 -43
rect 386 -44 387 -43
rect 387 -44 388 -43
rect 388 -44 389 -43
rect 389 -44 390 -43
rect 390 -44 391 -43
rect 391 -44 392 -43
rect 392 -44 393 -43
rect 393 -44 394 -43
rect 394 -44 395 -43
rect 395 -44 396 -43
rect 396 -44 397 -43
rect 397 -44 398 -43
rect 398 -44 399 -43
rect 399 -44 400 -43
rect 400 -44 401 -43
rect 401 -44 402 -43
rect 402 -44 403 -43
rect 403 -44 404 -43
rect 404 -44 405 -43
rect 405 -44 406 -43
rect 406 -44 407 -43
rect 407 -44 408 -43
rect 408 -44 409 -43
rect 409 -44 410 -43
rect 410 -44 411 -43
rect 411 -44 412 -43
rect 412 -44 413 -43
rect 413 -44 414 -43
rect 414 -44 415 -43
rect 415 -44 416 -43
rect 416 -44 417 -43
rect 417 -44 418 -43
rect 418 -44 419 -43
rect 419 -44 420 -43
rect 420 -44 421 -43
rect 421 -44 422 -43
rect 422 -44 423 -43
rect 423 -44 424 -43
rect 424 -44 425 -43
rect 425 -44 426 -43
rect 426 -44 427 -43
rect 427 -44 428 -43
rect 428 -44 429 -43
rect 429 -44 430 -43
rect 430 -44 431 -43
rect 431 -44 432 -43
rect 432 -44 433 -43
rect 433 -44 434 -43
rect 434 -44 435 -43
rect 435 -44 436 -43
rect 436 -44 437 -43
rect 437 -44 438 -43
rect 438 -44 439 -43
rect 439 -44 440 -43
rect 440 -44 441 -43
rect 441 -44 442 -43
rect 442 -44 443 -43
rect 443 -44 444 -43
rect 444 -44 445 -43
rect 445 -44 446 -43
rect 446 -44 447 -43
rect 447 -44 448 -43
rect 448 -44 449 -43
rect 449 -44 450 -43
rect 450 -44 451 -43
rect 451 -44 452 -43
rect 452 -44 453 -43
rect 453 -44 454 -43
rect 454 -44 455 -43
rect 455 -44 456 -43
rect 456 -44 457 -43
rect 457 -44 458 -43
rect 458 -44 459 -43
rect 459 -44 460 -43
rect 460 -44 461 -43
rect 461 -44 462 -43
rect 462 -44 463 -43
rect 463 -44 464 -43
rect 464 -44 465 -43
rect 465 -44 466 -43
rect 466 -44 467 -43
rect 467 -44 468 -43
rect 468 -44 469 -43
rect 469 -44 470 -43
rect 470 -44 471 -43
rect 471 -44 472 -43
rect 472 -44 473 -43
rect 473 -44 474 -43
rect 474 -44 475 -43
rect 475 -44 476 -43
rect 476 -44 477 -43
rect 477 -44 478 -43
rect 478 -44 479 -43
rect 479 -44 480 -43
rect 2 -45 3 -44
rect 3 -45 4 -44
rect 4 -45 5 -44
rect 5 -45 6 -44
rect 6 -45 7 -44
rect 7 -45 8 -44
rect 8 -45 9 -44
rect 9 -45 10 -44
rect 10 -45 11 -44
rect 11 -45 12 -44
rect 16 -45 17 -44
rect 22 -45 23 -44
rect 23 -45 24 -44
rect 24 -45 25 -44
rect 25 -45 26 -44
rect 26 -45 27 -44
rect 27 -45 28 -44
rect 28 -45 29 -44
rect 29 -45 30 -44
rect 30 -45 31 -44
rect 31 -45 32 -44
rect 32 -45 33 -44
rect 33 -45 34 -44
rect 34 -45 35 -44
rect 35 -45 36 -44
rect 36 -45 37 -44
rect 37 -45 38 -44
rect 38 -45 39 -44
rect 39 -45 40 -44
rect 40 -45 41 -44
rect 41 -45 42 -44
rect 42 -45 43 -44
rect 43 -45 44 -44
rect 48 -45 49 -44
rect 54 -45 55 -44
rect 55 -45 56 -44
rect 56 -45 57 -44
rect 57 -45 58 -44
rect 58 -45 59 -44
rect 59 -45 60 -44
rect 60 -45 61 -44
rect 61 -45 62 -44
rect 62 -45 63 -44
rect 63 -45 64 -44
rect 64 -45 65 -44
rect 65 -45 66 -44
rect 66 -45 67 -44
rect 67 -45 68 -44
rect 68 -45 69 -44
rect 69 -45 70 -44
rect 70 -45 71 -44
rect 71 -45 72 -44
rect 72 -45 73 -44
rect 73 -45 74 -44
rect 74 -45 75 -44
rect 75 -45 76 -44
rect 80 -45 81 -44
rect 86 -45 87 -44
rect 87 -45 88 -44
rect 88 -45 89 -44
rect 89 -45 90 -44
rect 90 -45 91 -44
rect 91 -45 92 -44
rect 92 -45 93 -44
rect 93 -45 94 -44
rect 94 -45 95 -44
rect 95 -45 96 -44
rect 96 -45 97 -44
rect 97 -45 98 -44
rect 98 -45 99 -44
rect 99 -45 100 -44
rect 100 -45 101 -44
rect 101 -45 102 -44
rect 102 -45 103 -44
rect 103 -45 104 -44
rect 104 -45 105 -44
rect 105 -45 106 -44
rect 106 -45 107 -44
rect 107 -45 108 -44
rect 112 -45 113 -44
rect 118 -45 119 -44
rect 119 -45 120 -44
rect 120 -45 121 -44
rect 121 -45 122 -44
rect 122 -45 123 -44
rect 123 -45 124 -44
rect 124 -45 125 -44
rect 125 -45 126 -44
rect 126 -45 127 -44
rect 127 -45 128 -44
rect 128 -45 129 -44
rect 129 -45 130 -44
rect 130 -45 131 -44
rect 131 -45 132 -44
rect 132 -45 133 -44
rect 133 -45 134 -44
rect 134 -45 135 -44
rect 135 -45 136 -44
rect 136 -45 137 -44
rect 137 -45 138 -44
rect 138 -45 139 -44
rect 139 -45 140 -44
rect 144 -45 145 -44
rect 150 -45 151 -44
rect 151 -45 152 -44
rect 152 -45 153 -44
rect 153 -45 154 -44
rect 154 -45 155 -44
rect 155 -45 156 -44
rect 156 -45 157 -44
rect 157 -45 158 -44
rect 158 -45 159 -44
rect 159 -45 160 -44
rect 160 -45 161 -44
rect 161 -45 162 -44
rect 162 -45 163 -44
rect 163 -45 164 -44
rect 164 -45 165 -44
rect 165 -45 166 -44
rect 166 -45 167 -44
rect 167 -45 168 -44
rect 168 -45 169 -44
rect 169 -45 170 -44
rect 170 -45 171 -44
rect 171 -45 172 -44
rect 176 -45 177 -44
rect 182 -45 183 -44
rect 183 -45 184 -44
rect 184 -45 185 -44
rect 185 -45 186 -44
rect 186 -45 187 -44
rect 187 -45 188 -44
rect 188 -45 189 -44
rect 189 -45 190 -44
rect 190 -45 191 -44
rect 191 -45 192 -44
rect 192 -45 193 -44
rect 193 -45 194 -44
rect 194 -45 195 -44
rect 195 -45 196 -44
rect 196 -45 197 -44
rect 197 -45 198 -44
rect 198 -45 199 -44
rect 199 -45 200 -44
rect 200 -45 201 -44
rect 201 -45 202 -44
rect 202 -45 203 -44
rect 203 -45 204 -44
rect 204 -45 205 -44
rect 205 -45 206 -44
rect 206 -45 207 -44
rect 207 -45 208 -44
rect 208 -45 209 -44
rect 209 -45 210 -44
rect 210 -45 211 -44
rect 211 -45 212 -44
rect 212 -45 213 -44
rect 213 -45 214 -44
rect 214 -45 215 -44
rect 215 -45 216 -44
rect 216 -45 217 -44
rect 217 -45 218 -44
rect 218 -45 219 -44
rect 219 -45 220 -44
rect 220 -45 221 -44
rect 221 -45 222 -44
rect 222 -45 223 -44
rect 223 -45 224 -44
rect 224 -45 225 -44
rect 225 -45 226 -44
rect 226 -45 227 -44
rect 227 -45 228 -44
rect 228 -45 229 -44
rect 229 -45 230 -44
rect 230 -45 231 -44
rect 231 -45 232 -44
rect 232 -45 233 -44
rect 233 -45 234 -44
rect 234 -45 235 -44
rect 235 -45 236 -44
rect 236 -45 237 -44
rect 237 -45 238 -44
rect 238 -45 239 -44
rect 239 -45 240 -44
rect 240 -45 241 -44
rect 241 -45 242 -44
rect 242 -45 243 -44
rect 243 -45 244 -44
rect 244 -45 245 -44
rect 245 -45 246 -44
rect 246 -45 247 -44
rect 247 -45 248 -44
rect 248 -45 249 -44
rect 249 -45 250 -44
rect 250 -45 251 -44
rect 251 -45 252 -44
rect 252 -45 253 -44
rect 253 -45 254 -44
rect 254 -45 255 -44
rect 255 -45 256 -44
rect 256 -45 257 -44
rect 257 -45 258 -44
rect 258 -45 259 -44
rect 259 -45 260 -44
rect 260 -45 261 -44
rect 261 -45 262 -44
rect 262 -45 263 -44
rect 263 -45 264 -44
rect 264 -45 265 -44
rect 265 -45 266 -44
rect 266 -45 267 -44
rect 267 -45 268 -44
rect 268 -45 269 -44
rect 269 -45 270 -44
rect 270 -45 271 -44
rect 271 -45 272 -44
rect 272 -45 273 -44
rect 273 -45 274 -44
rect 274 -45 275 -44
rect 275 -45 276 -44
rect 276 -45 277 -44
rect 277 -45 278 -44
rect 278 -45 279 -44
rect 279 -45 280 -44
rect 280 -45 281 -44
rect 281 -45 282 -44
rect 282 -45 283 -44
rect 283 -45 284 -44
rect 284 -45 285 -44
rect 285 -45 286 -44
rect 286 -45 287 -44
rect 287 -45 288 -44
rect 288 -45 289 -44
rect 289 -45 290 -44
rect 290 -45 291 -44
rect 291 -45 292 -44
rect 292 -45 293 -44
rect 293 -45 294 -44
rect 294 -45 295 -44
rect 295 -45 296 -44
rect 296 -45 297 -44
rect 297 -45 298 -44
rect 298 -45 299 -44
rect 299 -45 300 -44
rect 300 -45 301 -44
rect 301 -45 302 -44
rect 302 -45 303 -44
rect 303 -45 304 -44
rect 304 -45 305 -44
rect 305 -45 306 -44
rect 306 -45 307 -44
rect 307 -45 308 -44
rect 308 -45 309 -44
rect 309 -45 310 -44
rect 310 -45 311 -44
rect 311 -45 312 -44
rect 312 -45 313 -44
rect 313 -45 314 -44
rect 314 -45 315 -44
rect 315 -45 316 -44
rect 316 -45 317 -44
rect 317 -45 318 -44
rect 318 -45 319 -44
rect 319 -45 320 -44
rect 320 -45 321 -44
rect 321 -45 322 -44
rect 322 -45 323 -44
rect 323 -45 324 -44
rect 324 -45 325 -44
rect 325 -45 326 -44
rect 326 -45 327 -44
rect 327 -45 328 -44
rect 328 -45 329 -44
rect 329 -45 330 -44
rect 330 -45 331 -44
rect 331 -45 332 -44
rect 332 -45 333 -44
rect 333 -45 334 -44
rect 334 -45 335 -44
rect 335 -45 336 -44
rect 336 -45 337 -44
rect 337 -45 338 -44
rect 338 -45 339 -44
rect 339 -45 340 -44
rect 340 -45 341 -44
rect 341 -45 342 -44
rect 342 -45 343 -44
rect 343 -45 344 -44
rect 344 -45 345 -44
rect 345 -45 346 -44
rect 346 -45 347 -44
rect 347 -45 348 -44
rect 348 -45 349 -44
rect 349 -45 350 -44
rect 350 -45 351 -44
rect 351 -45 352 -44
rect 352 -45 353 -44
rect 353 -45 354 -44
rect 354 -45 355 -44
rect 355 -45 356 -44
rect 356 -45 357 -44
rect 357 -45 358 -44
rect 358 -45 359 -44
rect 359 -45 360 -44
rect 360 -45 361 -44
rect 361 -45 362 -44
rect 362 -45 363 -44
rect 363 -45 364 -44
rect 364 -45 365 -44
rect 365 -45 366 -44
rect 366 -45 367 -44
rect 367 -45 368 -44
rect 368 -45 369 -44
rect 369 -45 370 -44
rect 370 -45 371 -44
rect 371 -45 372 -44
rect 372 -45 373 -44
rect 373 -45 374 -44
rect 374 -45 375 -44
rect 375 -45 376 -44
rect 376 -45 377 -44
rect 377 -45 378 -44
rect 378 -45 379 -44
rect 379 -45 380 -44
rect 380 -45 381 -44
rect 381 -45 382 -44
rect 382 -45 383 -44
rect 383 -45 384 -44
rect 384 -45 385 -44
rect 385 -45 386 -44
rect 386 -45 387 -44
rect 387 -45 388 -44
rect 388 -45 389 -44
rect 389 -45 390 -44
rect 390 -45 391 -44
rect 391 -45 392 -44
rect 392 -45 393 -44
rect 393 -45 394 -44
rect 394 -45 395 -44
rect 395 -45 396 -44
rect 396 -45 397 -44
rect 397 -45 398 -44
rect 398 -45 399 -44
rect 399 -45 400 -44
rect 400 -45 401 -44
rect 401 -45 402 -44
rect 402 -45 403 -44
rect 403 -45 404 -44
rect 404 -45 405 -44
rect 405 -45 406 -44
rect 406 -45 407 -44
rect 407 -45 408 -44
rect 408 -45 409 -44
rect 409 -45 410 -44
rect 410 -45 411 -44
rect 411 -45 412 -44
rect 412 -45 413 -44
rect 413 -45 414 -44
rect 414 -45 415 -44
rect 415 -45 416 -44
rect 416 -45 417 -44
rect 417 -45 418 -44
rect 418 -45 419 -44
rect 419 -45 420 -44
rect 420 -45 421 -44
rect 421 -45 422 -44
rect 422 -45 423 -44
rect 423 -45 424 -44
rect 424 -45 425 -44
rect 425 -45 426 -44
rect 426 -45 427 -44
rect 427 -45 428 -44
rect 428 -45 429 -44
rect 429 -45 430 -44
rect 430 -45 431 -44
rect 431 -45 432 -44
rect 432 -45 433 -44
rect 433 -45 434 -44
rect 434 -45 435 -44
rect 435 -45 436 -44
rect 436 -45 437 -44
rect 437 -45 438 -44
rect 438 -45 439 -44
rect 439 -45 440 -44
rect 440 -45 441 -44
rect 441 -45 442 -44
rect 442 -45 443 -44
rect 443 -45 444 -44
rect 444 -45 445 -44
rect 445 -45 446 -44
rect 446 -45 447 -44
rect 447 -45 448 -44
rect 448 -45 449 -44
rect 449 -45 450 -44
rect 450 -45 451 -44
rect 451 -45 452 -44
rect 452 -45 453 -44
rect 453 -45 454 -44
rect 454 -45 455 -44
rect 455 -45 456 -44
rect 456 -45 457 -44
rect 457 -45 458 -44
rect 458 -45 459 -44
rect 459 -45 460 -44
rect 460 -45 461 -44
rect 461 -45 462 -44
rect 462 -45 463 -44
rect 463 -45 464 -44
rect 464 -45 465 -44
rect 465 -45 466 -44
rect 466 -45 467 -44
rect 467 -45 468 -44
rect 468 -45 469 -44
rect 469 -45 470 -44
rect 470 -45 471 -44
rect 471 -45 472 -44
rect 472 -45 473 -44
rect 473 -45 474 -44
rect 474 -45 475 -44
rect 475 -45 476 -44
rect 476 -45 477 -44
rect 477 -45 478 -44
rect 478 -45 479 -44
rect 479 -45 480 -44
rect 2 -46 3 -45
rect 3 -46 4 -45
rect 4 -46 5 -45
rect 5 -46 6 -45
rect 6 -46 7 -45
rect 7 -46 8 -45
rect 8 -46 9 -45
rect 9 -46 10 -45
rect 10 -46 11 -45
rect 15 -46 16 -45
rect 16 -46 17 -45
rect 17 -46 18 -45
rect 18 -46 19 -45
rect 22 -46 23 -45
rect 23 -46 24 -45
rect 24 -46 25 -45
rect 25 -46 26 -45
rect 26 -46 27 -45
rect 27 -46 28 -45
rect 28 -46 29 -45
rect 29 -46 30 -45
rect 30 -46 31 -45
rect 31 -46 32 -45
rect 32 -46 33 -45
rect 33 -46 34 -45
rect 34 -46 35 -45
rect 35 -46 36 -45
rect 36 -46 37 -45
rect 37 -46 38 -45
rect 38 -46 39 -45
rect 39 -46 40 -45
rect 40 -46 41 -45
rect 41 -46 42 -45
rect 42 -46 43 -45
rect 47 -46 48 -45
rect 48 -46 49 -45
rect 49 -46 50 -45
rect 50 -46 51 -45
rect 54 -46 55 -45
rect 55 -46 56 -45
rect 56 -46 57 -45
rect 57 -46 58 -45
rect 58 -46 59 -45
rect 59 -46 60 -45
rect 60 -46 61 -45
rect 61 -46 62 -45
rect 62 -46 63 -45
rect 63 -46 64 -45
rect 64 -46 65 -45
rect 65 -46 66 -45
rect 66 -46 67 -45
rect 67 -46 68 -45
rect 68 -46 69 -45
rect 69 -46 70 -45
rect 70 -46 71 -45
rect 71 -46 72 -45
rect 72 -46 73 -45
rect 73 -46 74 -45
rect 74 -46 75 -45
rect 79 -46 80 -45
rect 80 -46 81 -45
rect 81 -46 82 -45
rect 82 -46 83 -45
rect 86 -46 87 -45
rect 87 -46 88 -45
rect 88 -46 89 -45
rect 89 -46 90 -45
rect 90 -46 91 -45
rect 91 -46 92 -45
rect 92 -46 93 -45
rect 93 -46 94 -45
rect 94 -46 95 -45
rect 95 -46 96 -45
rect 96 -46 97 -45
rect 97 -46 98 -45
rect 98 -46 99 -45
rect 99 -46 100 -45
rect 100 -46 101 -45
rect 101 -46 102 -45
rect 102 -46 103 -45
rect 103 -46 104 -45
rect 104 -46 105 -45
rect 105 -46 106 -45
rect 106 -46 107 -45
rect 111 -46 112 -45
rect 112 -46 113 -45
rect 113 -46 114 -45
rect 114 -46 115 -45
rect 118 -46 119 -45
rect 119 -46 120 -45
rect 120 -46 121 -45
rect 121 -46 122 -45
rect 122 -46 123 -45
rect 123 -46 124 -45
rect 124 -46 125 -45
rect 125 -46 126 -45
rect 126 -46 127 -45
rect 127 -46 128 -45
rect 128 -46 129 -45
rect 129 -46 130 -45
rect 130 -46 131 -45
rect 131 -46 132 -45
rect 132 -46 133 -45
rect 133 -46 134 -45
rect 134 -46 135 -45
rect 135 -46 136 -45
rect 136 -46 137 -45
rect 137 -46 138 -45
rect 138 -46 139 -45
rect 143 -46 144 -45
rect 144 -46 145 -45
rect 145 -46 146 -45
rect 146 -46 147 -45
rect 150 -46 151 -45
rect 151 -46 152 -45
rect 152 -46 153 -45
rect 153 -46 154 -45
rect 154 -46 155 -45
rect 155 -46 156 -45
rect 156 -46 157 -45
rect 157 -46 158 -45
rect 158 -46 159 -45
rect 159 -46 160 -45
rect 160 -46 161 -45
rect 161 -46 162 -45
rect 162 -46 163 -45
rect 163 -46 164 -45
rect 164 -46 165 -45
rect 165 -46 166 -45
rect 166 -46 167 -45
rect 167 -46 168 -45
rect 168 -46 169 -45
rect 169 -46 170 -45
rect 170 -46 171 -45
rect 175 -46 176 -45
rect 176 -46 177 -45
rect 177 -46 178 -45
rect 178 -46 179 -45
rect 182 -46 183 -45
rect 183 -46 184 -45
rect 184 -46 185 -45
rect 185 -46 186 -45
rect 186 -46 187 -45
rect 187 -46 188 -45
rect 188 -46 189 -45
rect 189 -46 190 -45
rect 190 -46 191 -45
rect 191 -46 192 -45
rect 192 -46 193 -45
rect 193 -46 194 -45
rect 194 -46 195 -45
rect 195 -46 196 -45
rect 196 -46 197 -45
rect 197 -46 198 -45
rect 198 -46 199 -45
rect 199 -46 200 -45
rect 200 -46 201 -45
rect 201 -46 202 -45
rect 202 -46 203 -45
rect 203 -46 204 -45
rect 204 -46 205 -45
rect 205 -46 206 -45
rect 206 -46 207 -45
rect 207 -46 208 -45
rect 208 -46 209 -45
rect 209 -46 210 -45
rect 210 -46 211 -45
rect 211 -46 212 -45
rect 212 -46 213 -45
rect 213 -46 214 -45
rect 214 -46 215 -45
rect 215 -46 216 -45
rect 216 -46 217 -45
rect 217 -46 218 -45
rect 218 -46 219 -45
rect 219 -46 220 -45
rect 220 -46 221 -45
rect 221 -46 222 -45
rect 222 -46 223 -45
rect 223 -46 224 -45
rect 224 -46 225 -45
rect 225 -46 226 -45
rect 226 -46 227 -45
rect 227 -46 228 -45
rect 228 -46 229 -45
rect 229 -46 230 -45
rect 230 -46 231 -45
rect 231 -46 232 -45
rect 232 -46 233 -45
rect 233 -46 234 -45
rect 234 -46 235 -45
rect 235 -46 236 -45
rect 236 -46 237 -45
rect 237 -46 238 -45
rect 238 -46 239 -45
rect 239 -46 240 -45
rect 240 -46 241 -45
rect 241 -46 242 -45
rect 242 -46 243 -45
rect 243 -46 244 -45
rect 244 -46 245 -45
rect 245 -46 246 -45
rect 246 -46 247 -45
rect 247 -46 248 -45
rect 248 -46 249 -45
rect 249 -46 250 -45
rect 250 -46 251 -45
rect 251 -46 252 -45
rect 252 -46 253 -45
rect 253 -46 254 -45
rect 254 -46 255 -45
rect 255 -46 256 -45
rect 256 -46 257 -45
rect 257 -46 258 -45
rect 258 -46 259 -45
rect 259 -46 260 -45
rect 260 -46 261 -45
rect 261 -46 262 -45
rect 262 -46 263 -45
rect 263 -46 264 -45
rect 264 -46 265 -45
rect 265 -46 266 -45
rect 266 -46 267 -45
rect 267 -46 268 -45
rect 268 -46 269 -45
rect 269 -46 270 -45
rect 270 -46 271 -45
rect 271 -46 272 -45
rect 272 -46 273 -45
rect 273 -46 274 -45
rect 274 -46 275 -45
rect 275 -46 276 -45
rect 276 -46 277 -45
rect 277 -46 278 -45
rect 278 -46 279 -45
rect 279 -46 280 -45
rect 280 -46 281 -45
rect 281 -46 282 -45
rect 282 -46 283 -45
rect 283 -46 284 -45
rect 284 -46 285 -45
rect 285 -46 286 -45
rect 286 -46 287 -45
rect 287 -46 288 -45
rect 288 -46 289 -45
rect 289 -46 290 -45
rect 290 -46 291 -45
rect 291 -46 292 -45
rect 292 -46 293 -45
rect 293 -46 294 -45
rect 294 -46 295 -45
rect 295 -46 296 -45
rect 296 -46 297 -45
rect 297 -46 298 -45
rect 298 -46 299 -45
rect 299 -46 300 -45
rect 300 -46 301 -45
rect 301 -46 302 -45
rect 302 -46 303 -45
rect 303 -46 304 -45
rect 304 -46 305 -45
rect 305 -46 306 -45
rect 306 -46 307 -45
rect 307 -46 308 -45
rect 308 -46 309 -45
rect 309 -46 310 -45
rect 310 -46 311 -45
rect 311 -46 312 -45
rect 312 -46 313 -45
rect 313 -46 314 -45
rect 314 -46 315 -45
rect 315 -46 316 -45
rect 316 -46 317 -45
rect 317 -46 318 -45
rect 318 -46 319 -45
rect 319 -46 320 -45
rect 320 -46 321 -45
rect 321 -46 322 -45
rect 322 -46 323 -45
rect 323 -46 324 -45
rect 324 -46 325 -45
rect 325 -46 326 -45
rect 326 -46 327 -45
rect 327 -46 328 -45
rect 328 -46 329 -45
rect 329 -46 330 -45
rect 330 -46 331 -45
rect 331 -46 332 -45
rect 332 -46 333 -45
rect 333 -46 334 -45
rect 334 -46 335 -45
rect 335 -46 336 -45
rect 336 -46 337 -45
rect 337 -46 338 -45
rect 338 -46 339 -45
rect 339 -46 340 -45
rect 340 -46 341 -45
rect 341 -46 342 -45
rect 342 -46 343 -45
rect 343 -46 344 -45
rect 344 -46 345 -45
rect 345 -46 346 -45
rect 346 -46 347 -45
rect 347 -46 348 -45
rect 348 -46 349 -45
rect 349 -46 350 -45
rect 350 -46 351 -45
rect 351 -46 352 -45
rect 352 -46 353 -45
rect 353 -46 354 -45
rect 354 -46 355 -45
rect 355 -46 356 -45
rect 356 -46 357 -45
rect 357 -46 358 -45
rect 358 -46 359 -45
rect 359 -46 360 -45
rect 360 -46 361 -45
rect 361 -46 362 -45
rect 362 -46 363 -45
rect 363 -46 364 -45
rect 364 -46 365 -45
rect 365 -46 366 -45
rect 366 -46 367 -45
rect 367 -46 368 -45
rect 368 -46 369 -45
rect 369 -46 370 -45
rect 370 -46 371 -45
rect 371 -46 372 -45
rect 372 -46 373 -45
rect 373 -46 374 -45
rect 374 -46 375 -45
rect 375 -46 376 -45
rect 376 -46 377 -45
rect 377 -46 378 -45
rect 378 -46 379 -45
rect 379 -46 380 -45
rect 380 -46 381 -45
rect 381 -46 382 -45
rect 382 -46 383 -45
rect 383 -46 384 -45
rect 384 -46 385 -45
rect 385 -46 386 -45
rect 386 -46 387 -45
rect 387 -46 388 -45
rect 388 -46 389 -45
rect 389 -46 390 -45
rect 390 -46 391 -45
rect 391 -46 392 -45
rect 392 -46 393 -45
rect 393 -46 394 -45
rect 394 -46 395 -45
rect 395 -46 396 -45
rect 396 -46 397 -45
rect 397 -46 398 -45
rect 398 -46 399 -45
rect 399 -46 400 -45
rect 400 -46 401 -45
rect 401 -46 402 -45
rect 402 -46 403 -45
rect 403 -46 404 -45
rect 404 -46 405 -45
rect 405 -46 406 -45
rect 406 -46 407 -45
rect 407 -46 408 -45
rect 408 -46 409 -45
rect 409 -46 410 -45
rect 410 -46 411 -45
rect 411 -46 412 -45
rect 412 -46 413 -45
rect 413 -46 414 -45
rect 414 -46 415 -45
rect 415 -46 416 -45
rect 416 -46 417 -45
rect 417 -46 418 -45
rect 418 -46 419 -45
rect 419 -46 420 -45
rect 420 -46 421 -45
rect 421 -46 422 -45
rect 422 -46 423 -45
rect 423 -46 424 -45
rect 424 -46 425 -45
rect 425 -46 426 -45
rect 426 -46 427 -45
rect 427 -46 428 -45
rect 428 -46 429 -45
rect 429 -46 430 -45
rect 430 -46 431 -45
rect 431 -46 432 -45
rect 432 -46 433 -45
rect 433 -46 434 -45
rect 434 -46 435 -45
rect 435 -46 436 -45
rect 436 -46 437 -45
rect 437 -46 438 -45
rect 438 -46 439 -45
rect 439 -46 440 -45
rect 440 -46 441 -45
rect 441 -46 442 -45
rect 442 -46 443 -45
rect 443 -46 444 -45
rect 444 -46 445 -45
rect 445 -46 446 -45
rect 446 -46 447 -45
rect 447 -46 448 -45
rect 448 -46 449 -45
rect 449 -46 450 -45
rect 450 -46 451 -45
rect 451 -46 452 -45
rect 452 -46 453 -45
rect 453 -46 454 -45
rect 454 -46 455 -45
rect 455 -46 456 -45
rect 456 -46 457 -45
rect 457 -46 458 -45
rect 458 -46 459 -45
rect 459 -46 460 -45
rect 460 -46 461 -45
rect 461 -46 462 -45
rect 462 -46 463 -45
rect 463 -46 464 -45
rect 464 -46 465 -45
rect 465 -46 466 -45
rect 466 -46 467 -45
rect 467 -46 468 -45
rect 468 -46 469 -45
rect 469 -46 470 -45
rect 470 -46 471 -45
rect 471 -46 472 -45
rect 472 -46 473 -45
rect 473 -46 474 -45
rect 474 -46 475 -45
rect 475 -46 476 -45
rect 476 -46 477 -45
rect 477 -46 478 -45
rect 478 -46 479 -45
rect 479 -46 480 -45
rect 2 -47 3 -46
rect 3 -47 4 -46
rect 4 -47 5 -46
rect 5 -47 6 -46
rect 6 -47 7 -46
rect 7 -47 8 -46
rect 8 -47 9 -46
rect 9 -47 10 -46
rect 10 -47 11 -46
rect 14 -47 15 -46
rect 15 -47 16 -46
rect 16 -47 17 -46
rect 17 -47 18 -46
rect 18 -47 19 -46
rect 19 -47 20 -46
rect 22 -47 23 -46
rect 23 -47 24 -46
rect 24 -47 25 -46
rect 25 -47 26 -46
rect 26 -47 27 -46
rect 27 -47 28 -46
rect 28 -47 29 -46
rect 29 -47 30 -46
rect 30 -47 31 -46
rect 34 -47 35 -46
rect 35 -47 36 -46
rect 36 -47 37 -46
rect 37 -47 38 -46
rect 38 -47 39 -46
rect 39 -47 40 -46
rect 40 -47 41 -46
rect 41 -47 42 -46
rect 42 -47 43 -46
rect 46 -47 47 -46
rect 47 -47 48 -46
rect 48 -47 49 -46
rect 49 -47 50 -46
rect 50 -47 51 -46
rect 51 -47 52 -46
rect 54 -47 55 -46
rect 55 -47 56 -46
rect 56 -47 57 -46
rect 57 -47 58 -46
rect 58 -47 59 -46
rect 59 -47 60 -46
rect 60 -47 61 -46
rect 61 -47 62 -46
rect 62 -47 63 -46
rect 66 -47 67 -46
rect 67 -47 68 -46
rect 68 -47 69 -46
rect 69 -47 70 -46
rect 70 -47 71 -46
rect 71 -47 72 -46
rect 72 -47 73 -46
rect 73 -47 74 -46
rect 74 -47 75 -46
rect 78 -47 79 -46
rect 79 -47 80 -46
rect 80 -47 81 -46
rect 81 -47 82 -46
rect 82 -47 83 -46
rect 83 -47 84 -46
rect 86 -47 87 -46
rect 87 -47 88 -46
rect 88 -47 89 -46
rect 89 -47 90 -46
rect 90 -47 91 -46
rect 91 -47 92 -46
rect 92 -47 93 -46
rect 93 -47 94 -46
rect 94 -47 95 -46
rect 98 -47 99 -46
rect 99 -47 100 -46
rect 100 -47 101 -46
rect 101 -47 102 -46
rect 102 -47 103 -46
rect 103 -47 104 -46
rect 104 -47 105 -46
rect 105 -47 106 -46
rect 106 -47 107 -46
rect 110 -47 111 -46
rect 111 -47 112 -46
rect 112 -47 113 -46
rect 113 -47 114 -46
rect 114 -47 115 -46
rect 115 -47 116 -46
rect 118 -47 119 -46
rect 119 -47 120 -46
rect 120 -47 121 -46
rect 121 -47 122 -46
rect 122 -47 123 -46
rect 123 -47 124 -46
rect 124 -47 125 -46
rect 125 -47 126 -46
rect 126 -47 127 -46
rect 130 -47 131 -46
rect 131 -47 132 -46
rect 132 -47 133 -46
rect 133 -47 134 -46
rect 134 -47 135 -46
rect 135 -47 136 -46
rect 136 -47 137 -46
rect 137 -47 138 -46
rect 138 -47 139 -46
rect 142 -47 143 -46
rect 143 -47 144 -46
rect 144 -47 145 -46
rect 145 -47 146 -46
rect 146 -47 147 -46
rect 147 -47 148 -46
rect 150 -47 151 -46
rect 151 -47 152 -46
rect 152 -47 153 -46
rect 153 -47 154 -46
rect 154 -47 155 -46
rect 155 -47 156 -46
rect 156 -47 157 -46
rect 157 -47 158 -46
rect 158 -47 159 -46
rect 162 -47 163 -46
rect 163 -47 164 -46
rect 164 -47 165 -46
rect 165 -47 166 -46
rect 166 -47 167 -46
rect 167 -47 168 -46
rect 168 -47 169 -46
rect 169 -47 170 -46
rect 170 -47 171 -46
rect 174 -47 175 -46
rect 175 -47 176 -46
rect 176 -47 177 -46
rect 177 -47 178 -46
rect 178 -47 179 -46
rect 179 -47 180 -46
rect 182 -47 183 -46
rect 183 -47 184 -46
rect 184 -47 185 -46
rect 185 -47 186 -46
rect 186 -47 187 -46
rect 187 -47 188 -46
rect 188 -47 189 -46
rect 189 -47 190 -46
rect 190 -47 191 -46
rect 191 -47 192 -46
rect 192 -47 193 -46
rect 193 -47 194 -46
rect 194 -47 195 -46
rect 195 -47 196 -46
rect 196 -47 197 -46
rect 197 -47 198 -46
rect 198 -47 199 -46
rect 199 -47 200 -46
rect 200 -47 201 -46
rect 201 -47 202 -46
rect 202 -47 203 -46
rect 203 -47 204 -46
rect 204 -47 205 -46
rect 205 -47 206 -46
rect 206 -47 207 -46
rect 207 -47 208 -46
rect 208 -47 209 -46
rect 209 -47 210 -46
rect 210 -47 211 -46
rect 211 -47 212 -46
rect 212 -47 213 -46
rect 213 -47 214 -46
rect 214 -47 215 -46
rect 215 -47 216 -46
rect 216 -47 217 -46
rect 217 -47 218 -46
rect 218 -47 219 -46
rect 219 -47 220 -46
rect 220 -47 221 -46
rect 221 -47 222 -46
rect 222 -47 223 -46
rect 223 -47 224 -46
rect 224 -47 225 -46
rect 225 -47 226 -46
rect 226 -47 227 -46
rect 227 -47 228 -46
rect 228 -47 229 -46
rect 229 -47 230 -46
rect 230 -47 231 -46
rect 231 -47 232 -46
rect 232 -47 233 -46
rect 233 -47 234 -46
rect 234 -47 235 -46
rect 235 -47 236 -46
rect 236 -47 237 -46
rect 237 -47 238 -46
rect 238 -47 239 -46
rect 239 -47 240 -46
rect 240 -47 241 -46
rect 241 -47 242 -46
rect 242 -47 243 -46
rect 243 -47 244 -46
rect 244 -47 245 -46
rect 245 -47 246 -46
rect 246 -47 247 -46
rect 247 -47 248 -46
rect 248 -47 249 -46
rect 249 -47 250 -46
rect 250 -47 251 -46
rect 251 -47 252 -46
rect 252 -47 253 -46
rect 253 -47 254 -46
rect 254 -47 255 -46
rect 255 -47 256 -46
rect 256 -47 257 -46
rect 257 -47 258 -46
rect 258 -47 259 -46
rect 259 -47 260 -46
rect 260 -47 261 -46
rect 261 -47 262 -46
rect 262 -47 263 -46
rect 263 -47 264 -46
rect 264 -47 265 -46
rect 265 -47 266 -46
rect 266 -47 267 -46
rect 267 -47 268 -46
rect 268 -47 269 -46
rect 269 -47 270 -46
rect 270 -47 271 -46
rect 271 -47 272 -46
rect 272 -47 273 -46
rect 273 -47 274 -46
rect 274 -47 275 -46
rect 275 -47 276 -46
rect 276 -47 277 -46
rect 277 -47 278 -46
rect 278 -47 279 -46
rect 279 -47 280 -46
rect 280 -47 281 -46
rect 281 -47 282 -46
rect 282 -47 283 -46
rect 283 -47 284 -46
rect 284 -47 285 -46
rect 285 -47 286 -46
rect 286 -47 287 -46
rect 287 -47 288 -46
rect 288 -47 289 -46
rect 289 -47 290 -46
rect 290 -47 291 -46
rect 291 -47 292 -46
rect 292 -47 293 -46
rect 293 -47 294 -46
rect 294 -47 295 -46
rect 295 -47 296 -46
rect 296 -47 297 -46
rect 297 -47 298 -46
rect 298 -47 299 -46
rect 299 -47 300 -46
rect 300 -47 301 -46
rect 301 -47 302 -46
rect 302 -47 303 -46
rect 303 -47 304 -46
rect 304 -47 305 -46
rect 305 -47 306 -46
rect 306 -47 307 -46
rect 307 -47 308 -46
rect 308 -47 309 -46
rect 309 -47 310 -46
rect 310 -47 311 -46
rect 311 -47 312 -46
rect 312 -47 313 -46
rect 313 -47 314 -46
rect 314 -47 315 -46
rect 315 -47 316 -46
rect 316 -47 317 -46
rect 317 -47 318 -46
rect 318 -47 319 -46
rect 319 -47 320 -46
rect 320 -47 321 -46
rect 321 -47 322 -46
rect 322 -47 323 -46
rect 323 -47 324 -46
rect 324 -47 325 -46
rect 325 -47 326 -46
rect 326 -47 327 -46
rect 327 -47 328 -46
rect 328 -47 329 -46
rect 329 -47 330 -46
rect 330 -47 331 -46
rect 331 -47 332 -46
rect 332 -47 333 -46
rect 333 -47 334 -46
rect 334 -47 335 -46
rect 335 -47 336 -46
rect 336 -47 337 -46
rect 337 -47 338 -46
rect 338 -47 339 -46
rect 339 -47 340 -46
rect 340 -47 341 -46
rect 341 -47 342 -46
rect 342 -47 343 -46
rect 343 -47 344 -46
rect 344 -47 345 -46
rect 345 -47 346 -46
rect 346 -47 347 -46
rect 347 -47 348 -46
rect 348 -47 349 -46
rect 349 -47 350 -46
rect 350 -47 351 -46
rect 351 -47 352 -46
rect 352 -47 353 -46
rect 353 -47 354 -46
rect 354 -47 355 -46
rect 355 -47 356 -46
rect 356 -47 357 -46
rect 357 -47 358 -46
rect 358 -47 359 -46
rect 359 -47 360 -46
rect 360 -47 361 -46
rect 361 -47 362 -46
rect 362 -47 363 -46
rect 363 -47 364 -46
rect 364 -47 365 -46
rect 365 -47 366 -46
rect 366 -47 367 -46
rect 367 -47 368 -46
rect 368 -47 369 -46
rect 369 -47 370 -46
rect 370 -47 371 -46
rect 371 -47 372 -46
rect 372 -47 373 -46
rect 373 -47 374 -46
rect 374 -47 375 -46
rect 375 -47 376 -46
rect 376 -47 377 -46
rect 377 -47 378 -46
rect 378 -47 379 -46
rect 379 -47 380 -46
rect 380 -47 381 -46
rect 381 -47 382 -46
rect 382 -47 383 -46
rect 383 -47 384 -46
rect 384 -47 385 -46
rect 385 -47 386 -46
rect 386 -47 387 -46
rect 387 -47 388 -46
rect 388 -47 389 -46
rect 389 -47 390 -46
rect 390 -47 391 -46
rect 391 -47 392 -46
rect 392 -47 393 -46
rect 393 -47 394 -46
rect 394 -47 395 -46
rect 395 -47 396 -46
rect 396 -47 397 -46
rect 397 -47 398 -46
rect 398 -47 399 -46
rect 399 -47 400 -46
rect 400 -47 401 -46
rect 401 -47 402 -46
rect 402 -47 403 -46
rect 403 -47 404 -46
rect 404 -47 405 -46
rect 405 -47 406 -46
rect 406 -47 407 -46
rect 407 -47 408 -46
rect 408 -47 409 -46
rect 409 -47 410 -46
rect 410 -47 411 -46
rect 411 -47 412 -46
rect 412 -47 413 -46
rect 413 -47 414 -46
rect 414 -47 415 -46
rect 415 -47 416 -46
rect 416 -47 417 -46
rect 417 -47 418 -46
rect 418 -47 419 -46
rect 419 -47 420 -46
rect 420 -47 421 -46
rect 421 -47 422 -46
rect 422 -47 423 -46
rect 423 -47 424 -46
rect 424 -47 425 -46
rect 425 -47 426 -46
rect 426 -47 427 -46
rect 427 -47 428 -46
rect 428 -47 429 -46
rect 429 -47 430 -46
rect 430 -47 431 -46
rect 431 -47 432 -46
rect 432 -47 433 -46
rect 433 -47 434 -46
rect 434 -47 435 -46
rect 435 -47 436 -46
rect 436 -47 437 -46
rect 437 -47 438 -46
rect 438 -47 439 -46
rect 439 -47 440 -46
rect 440 -47 441 -46
rect 441 -47 442 -46
rect 442 -47 443 -46
rect 443 -47 444 -46
rect 444 -47 445 -46
rect 445 -47 446 -46
rect 446 -47 447 -46
rect 447 -47 448 -46
rect 448 -47 449 -46
rect 449 -47 450 -46
rect 450 -47 451 -46
rect 451 -47 452 -46
rect 452 -47 453 -46
rect 453 -47 454 -46
rect 454 -47 455 -46
rect 455 -47 456 -46
rect 456 -47 457 -46
rect 457 -47 458 -46
rect 458 -47 459 -46
rect 459 -47 460 -46
rect 460 -47 461 -46
rect 461 -47 462 -46
rect 462 -47 463 -46
rect 463 -47 464 -46
rect 464 -47 465 -46
rect 465 -47 466 -46
rect 466 -47 467 -46
rect 467 -47 468 -46
rect 468 -47 469 -46
rect 469 -47 470 -46
rect 470 -47 471 -46
rect 471 -47 472 -46
rect 472 -47 473 -46
rect 473 -47 474 -46
rect 474 -47 475 -46
rect 475 -47 476 -46
rect 476 -47 477 -46
rect 477 -47 478 -46
rect 478 -47 479 -46
rect 479 -47 480 -46
rect 2 -48 3 -47
rect 3 -48 4 -47
rect 4 -48 5 -47
rect 5 -48 6 -47
rect 6 -48 7 -47
rect 7 -48 8 -47
rect 8 -48 9 -47
rect 9 -48 10 -47
rect 10 -48 11 -47
rect 11 -48 12 -47
rect 12 -48 13 -47
rect 13 -48 14 -47
rect 14 -48 15 -47
rect 15 -48 16 -47
rect 16 -48 17 -47
rect 17 -48 18 -47
rect 18 -48 19 -47
rect 19 -48 20 -47
rect 20 -48 21 -47
rect 21 -48 22 -47
rect 22 -48 23 -47
rect 23 -48 24 -47
rect 24 -48 25 -47
rect 25 -48 26 -47
rect 26 -48 27 -47
rect 27 -48 28 -47
rect 28 -48 29 -47
rect 29 -48 30 -47
rect 30 -48 31 -47
rect 34 -48 35 -47
rect 35 -48 36 -47
rect 36 -48 37 -47
rect 37 -48 38 -47
rect 38 -48 39 -47
rect 39 -48 40 -47
rect 40 -48 41 -47
rect 41 -48 42 -47
rect 42 -48 43 -47
rect 43 -48 44 -47
rect 44 -48 45 -47
rect 45 -48 46 -47
rect 46 -48 47 -47
rect 47 -48 48 -47
rect 48 -48 49 -47
rect 49 -48 50 -47
rect 50 -48 51 -47
rect 51 -48 52 -47
rect 52 -48 53 -47
rect 53 -48 54 -47
rect 54 -48 55 -47
rect 55 -48 56 -47
rect 56 -48 57 -47
rect 57 -48 58 -47
rect 58 -48 59 -47
rect 59 -48 60 -47
rect 60 -48 61 -47
rect 61 -48 62 -47
rect 62 -48 63 -47
rect 66 -48 67 -47
rect 67 -48 68 -47
rect 68 -48 69 -47
rect 69 -48 70 -47
rect 70 -48 71 -47
rect 71 -48 72 -47
rect 72 -48 73 -47
rect 73 -48 74 -47
rect 74 -48 75 -47
rect 75 -48 76 -47
rect 76 -48 77 -47
rect 77 -48 78 -47
rect 78 -48 79 -47
rect 79 -48 80 -47
rect 80 -48 81 -47
rect 81 -48 82 -47
rect 82 -48 83 -47
rect 83 -48 84 -47
rect 84 -48 85 -47
rect 85 -48 86 -47
rect 86 -48 87 -47
rect 87 -48 88 -47
rect 88 -48 89 -47
rect 89 -48 90 -47
rect 90 -48 91 -47
rect 91 -48 92 -47
rect 92 -48 93 -47
rect 93 -48 94 -47
rect 94 -48 95 -47
rect 98 -48 99 -47
rect 99 -48 100 -47
rect 100 -48 101 -47
rect 101 -48 102 -47
rect 102 -48 103 -47
rect 103 -48 104 -47
rect 104 -48 105 -47
rect 105 -48 106 -47
rect 106 -48 107 -47
rect 107 -48 108 -47
rect 108 -48 109 -47
rect 109 -48 110 -47
rect 110 -48 111 -47
rect 111 -48 112 -47
rect 112 -48 113 -47
rect 113 -48 114 -47
rect 114 -48 115 -47
rect 115 -48 116 -47
rect 116 -48 117 -47
rect 117 -48 118 -47
rect 118 -48 119 -47
rect 119 -48 120 -47
rect 120 -48 121 -47
rect 121 -48 122 -47
rect 122 -48 123 -47
rect 123 -48 124 -47
rect 124 -48 125 -47
rect 125 -48 126 -47
rect 126 -48 127 -47
rect 130 -48 131 -47
rect 131 -48 132 -47
rect 132 -48 133 -47
rect 133 -48 134 -47
rect 134 -48 135 -47
rect 135 -48 136 -47
rect 136 -48 137 -47
rect 137 -48 138 -47
rect 138 -48 139 -47
rect 139 -48 140 -47
rect 140 -48 141 -47
rect 141 -48 142 -47
rect 142 -48 143 -47
rect 143 -48 144 -47
rect 144 -48 145 -47
rect 145 -48 146 -47
rect 146 -48 147 -47
rect 147 -48 148 -47
rect 148 -48 149 -47
rect 149 -48 150 -47
rect 150 -48 151 -47
rect 151 -48 152 -47
rect 152 -48 153 -47
rect 153 -48 154 -47
rect 154 -48 155 -47
rect 155 -48 156 -47
rect 156 -48 157 -47
rect 157 -48 158 -47
rect 158 -48 159 -47
rect 162 -48 163 -47
rect 163 -48 164 -47
rect 164 -48 165 -47
rect 165 -48 166 -47
rect 166 -48 167 -47
rect 167 -48 168 -47
rect 168 -48 169 -47
rect 169 -48 170 -47
rect 170 -48 171 -47
rect 171 -48 172 -47
rect 172 -48 173 -47
rect 173 -48 174 -47
rect 174 -48 175 -47
rect 175 -48 176 -47
rect 176 -48 177 -47
rect 177 -48 178 -47
rect 178 -48 179 -47
rect 179 -48 180 -47
rect 180 -48 181 -47
rect 181 -48 182 -47
rect 182 -48 183 -47
rect 183 -48 184 -47
rect 184 -48 185 -47
rect 185 -48 186 -47
rect 186 -48 187 -47
rect 187 -48 188 -47
rect 188 -48 189 -47
rect 189 -48 190 -47
rect 190 -48 191 -47
rect 191 -48 192 -47
rect 192 -48 193 -47
rect 193 -48 194 -47
rect 194 -48 195 -47
rect 195 -48 196 -47
rect 196 -48 197 -47
rect 197 -48 198 -47
rect 198 -48 199 -47
rect 199 -48 200 -47
rect 200 -48 201 -47
rect 201 -48 202 -47
rect 202 -48 203 -47
rect 203 -48 204 -47
rect 204 -48 205 -47
rect 205 -48 206 -47
rect 206 -48 207 -47
rect 207 -48 208 -47
rect 208 -48 209 -47
rect 209 -48 210 -47
rect 210 -48 211 -47
rect 211 -48 212 -47
rect 212 -48 213 -47
rect 213 -48 214 -47
rect 214 -48 215 -47
rect 215 -48 216 -47
rect 216 -48 217 -47
rect 217 -48 218 -47
rect 218 -48 219 -47
rect 219 -48 220 -47
rect 220 -48 221 -47
rect 221 -48 222 -47
rect 222 -48 223 -47
rect 223 -48 224 -47
rect 224 -48 225 -47
rect 225 -48 226 -47
rect 226 -48 227 -47
rect 227 -48 228 -47
rect 228 -48 229 -47
rect 229 -48 230 -47
rect 230 -48 231 -47
rect 231 -48 232 -47
rect 232 -48 233 -47
rect 233 -48 234 -47
rect 234 -48 235 -47
rect 235 -48 236 -47
rect 236 -48 237 -47
rect 237 -48 238 -47
rect 238 -48 239 -47
rect 239 -48 240 -47
rect 240 -48 241 -47
rect 241 -48 242 -47
rect 242 -48 243 -47
rect 243 -48 244 -47
rect 244 -48 245 -47
rect 245 -48 246 -47
rect 246 -48 247 -47
rect 247 -48 248 -47
rect 248 -48 249 -47
rect 249 -48 250 -47
rect 250 -48 251 -47
rect 251 -48 252 -47
rect 252 -48 253 -47
rect 253 -48 254 -47
rect 254 -48 255 -47
rect 255 -48 256 -47
rect 256 -48 257 -47
rect 257 -48 258 -47
rect 258 -48 259 -47
rect 259 -48 260 -47
rect 260 -48 261 -47
rect 261 -48 262 -47
rect 262 -48 263 -47
rect 263 -48 264 -47
rect 264 -48 265 -47
rect 265 -48 266 -47
rect 266 -48 267 -47
rect 267 -48 268 -47
rect 268 -48 269 -47
rect 269 -48 270 -47
rect 270 -48 271 -47
rect 271 -48 272 -47
rect 272 -48 273 -47
rect 273 -48 274 -47
rect 274 -48 275 -47
rect 275 -48 276 -47
rect 276 -48 277 -47
rect 277 -48 278 -47
rect 278 -48 279 -47
rect 279 -48 280 -47
rect 280 -48 281 -47
rect 281 -48 282 -47
rect 282 -48 283 -47
rect 283 -48 284 -47
rect 284 -48 285 -47
rect 285 -48 286 -47
rect 286 -48 287 -47
rect 287 -48 288 -47
rect 288 -48 289 -47
rect 289 -48 290 -47
rect 290 -48 291 -47
rect 291 -48 292 -47
rect 292 -48 293 -47
rect 293 -48 294 -47
rect 294 -48 295 -47
rect 295 -48 296 -47
rect 296 -48 297 -47
rect 297 -48 298 -47
rect 298 -48 299 -47
rect 299 -48 300 -47
rect 300 -48 301 -47
rect 301 -48 302 -47
rect 302 -48 303 -47
rect 303 -48 304 -47
rect 304 -48 305 -47
rect 305 -48 306 -47
rect 306 -48 307 -47
rect 307 -48 308 -47
rect 308 -48 309 -47
rect 309 -48 310 -47
rect 310 -48 311 -47
rect 311 -48 312 -47
rect 312 -48 313 -47
rect 313 -48 314 -47
rect 314 -48 315 -47
rect 315 -48 316 -47
rect 316 -48 317 -47
rect 317 -48 318 -47
rect 318 -48 319 -47
rect 319 -48 320 -47
rect 320 -48 321 -47
rect 321 -48 322 -47
rect 322 -48 323 -47
rect 323 -48 324 -47
rect 324 -48 325 -47
rect 325 -48 326 -47
rect 326 -48 327 -47
rect 327 -48 328 -47
rect 328 -48 329 -47
rect 329 -48 330 -47
rect 330 -48 331 -47
rect 331 -48 332 -47
rect 332 -48 333 -47
rect 333 -48 334 -47
rect 334 -48 335 -47
rect 335 -48 336 -47
rect 336 -48 337 -47
rect 337 -48 338 -47
rect 338 -48 339 -47
rect 339 -48 340 -47
rect 340 -48 341 -47
rect 341 -48 342 -47
rect 342 -48 343 -47
rect 343 -48 344 -47
rect 344 -48 345 -47
rect 345 -48 346 -47
rect 346 -48 347 -47
rect 347 -48 348 -47
rect 348 -48 349 -47
rect 349 -48 350 -47
rect 350 -48 351 -47
rect 351 -48 352 -47
rect 352 -48 353 -47
rect 353 -48 354 -47
rect 354 -48 355 -47
rect 355 -48 356 -47
rect 356 -48 357 -47
rect 357 -48 358 -47
rect 358 -48 359 -47
rect 359 -48 360 -47
rect 360 -48 361 -47
rect 361 -48 362 -47
rect 362 -48 363 -47
rect 363 -48 364 -47
rect 364 -48 365 -47
rect 365 -48 366 -47
rect 366 -48 367 -47
rect 367 -48 368 -47
rect 368 -48 369 -47
rect 369 -48 370 -47
rect 370 -48 371 -47
rect 371 -48 372 -47
rect 372 -48 373 -47
rect 373 -48 374 -47
rect 374 -48 375 -47
rect 375 -48 376 -47
rect 376 -48 377 -47
rect 377 -48 378 -47
rect 378 -48 379 -47
rect 379 -48 380 -47
rect 380 -48 381 -47
rect 381 -48 382 -47
rect 382 -48 383 -47
rect 383 -48 384 -47
rect 384 -48 385 -47
rect 385 -48 386 -47
rect 386 -48 387 -47
rect 387 -48 388 -47
rect 388 -48 389 -47
rect 389 -48 390 -47
rect 390 -48 391 -47
rect 391 -48 392 -47
rect 392 -48 393 -47
rect 393 -48 394 -47
rect 394 -48 395 -47
rect 395 -48 396 -47
rect 396 -48 397 -47
rect 397 -48 398 -47
rect 398 -48 399 -47
rect 399 -48 400 -47
rect 400 -48 401 -47
rect 401 -48 402 -47
rect 402 -48 403 -47
rect 403 -48 404 -47
rect 404 -48 405 -47
rect 405 -48 406 -47
rect 406 -48 407 -47
rect 407 -48 408 -47
rect 408 -48 409 -47
rect 409 -48 410 -47
rect 410 -48 411 -47
rect 411 -48 412 -47
rect 412 -48 413 -47
rect 413 -48 414 -47
rect 414 -48 415 -47
rect 415 -48 416 -47
rect 416 -48 417 -47
rect 417 -48 418 -47
rect 418 -48 419 -47
rect 419 -48 420 -47
rect 420 -48 421 -47
rect 421 -48 422 -47
rect 422 -48 423 -47
rect 423 -48 424 -47
rect 424 -48 425 -47
rect 425 -48 426 -47
rect 426 -48 427 -47
rect 427 -48 428 -47
rect 428 -48 429 -47
rect 429 -48 430 -47
rect 430 -48 431 -47
rect 431 -48 432 -47
rect 432 -48 433 -47
rect 433 -48 434 -47
rect 434 -48 435 -47
rect 435 -48 436 -47
rect 436 -48 437 -47
rect 437 -48 438 -47
rect 438 -48 439 -47
rect 439 -48 440 -47
rect 440 -48 441 -47
rect 441 -48 442 -47
rect 442 -48 443 -47
rect 443 -48 444 -47
rect 444 -48 445 -47
rect 445 -48 446 -47
rect 446 -48 447 -47
rect 447 -48 448 -47
rect 448 -48 449 -47
rect 449 -48 450 -47
rect 450 -48 451 -47
rect 451 -48 452 -47
rect 452 -48 453 -47
rect 453 -48 454 -47
rect 454 -48 455 -47
rect 455 -48 456 -47
rect 456 -48 457 -47
rect 457 -48 458 -47
rect 458 -48 459 -47
rect 459 -48 460 -47
rect 460 -48 461 -47
rect 461 -48 462 -47
rect 462 -48 463 -47
rect 463 -48 464 -47
rect 464 -48 465 -47
rect 465 -48 466 -47
rect 466 -48 467 -47
rect 467 -48 468 -47
rect 468 -48 469 -47
rect 469 -48 470 -47
rect 470 -48 471 -47
rect 471 -48 472 -47
rect 472 -48 473 -47
rect 473 -48 474 -47
rect 474 -48 475 -47
rect 475 -48 476 -47
rect 476 -48 477 -47
rect 477 -48 478 -47
rect 478 -48 479 -47
rect 479 -48 480 -47
rect 2 -49 3 -48
rect 3 -49 4 -48
rect 4 -49 5 -48
rect 5 -49 6 -48
rect 6 -49 7 -48
rect 7 -49 8 -48
rect 8 -49 9 -48
rect 9 -49 10 -48
rect 10 -49 11 -48
rect 11 -49 12 -48
rect 12 -49 13 -48
rect 13 -49 14 -48
rect 14 -49 15 -48
rect 15 -49 16 -48
rect 16 -49 17 -48
rect 17 -49 18 -48
rect 18 -49 19 -48
rect 19 -49 20 -48
rect 20 -49 21 -48
rect 21 -49 22 -48
rect 22 -49 23 -48
rect 23 -49 24 -48
rect 24 -49 25 -48
rect 25 -49 26 -48
rect 26 -49 27 -48
rect 27 -49 28 -48
rect 28 -49 29 -48
rect 29 -49 30 -48
rect 30 -49 31 -48
rect 35 -49 36 -48
rect 36 -49 37 -48
rect 37 -49 38 -48
rect 38 -49 39 -48
rect 39 -49 40 -48
rect 40 -49 41 -48
rect 41 -49 42 -48
rect 42 -49 43 -48
rect 43 -49 44 -48
rect 44 -49 45 -48
rect 45 -49 46 -48
rect 46 -49 47 -48
rect 47 -49 48 -48
rect 48 -49 49 -48
rect 49 -49 50 -48
rect 50 -49 51 -48
rect 51 -49 52 -48
rect 52 -49 53 -48
rect 53 -49 54 -48
rect 54 -49 55 -48
rect 55 -49 56 -48
rect 56 -49 57 -48
rect 57 -49 58 -48
rect 58 -49 59 -48
rect 59 -49 60 -48
rect 60 -49 61 -48
rect 61 -49 62 -48
rect 62 -49 63 -48
rect 67 -49 68 -48
rect 68 -49 69 -48
rect 69 -49 70 -48
rect 70 -49 71 -48
rect 71 -49 72 -48
rect 72 -49 73 -48
rect 73 -49 74 -48
rect 74 -49 75 -48
rect 75 -49 76 -48
rect 76 -49 77 -48
rect 77 -49 78 -48
rect 78 -49 79 -48
rect 79 -49 80 -48
rect 80 -49 81 -48
rect 81 -49 82 -48
rect 82 -49 83 -48
rect 83 -49 84 -48
rect 84 -49 85 -48
rect 85 -49 86 -48
rect 86 -49 87 -48
rect 87 -49 88 -48
rect 88 -49 89 -48
rect 89 -49 90 -48
rect 90 -49 91 -48
rect 91 -49 92 -48
rect 92 -49 93 -48
rect 93 -49 94 -48
rect 94 -49 95 -48
rect 99 -49 100 -48
rect 100 -49 101 -48
rect 101 -49 102 -48
rect 102 -49 103 -48
rect 103 -49 104 -48
rect 104 -49 105 -48
rect 105 -49 106 -48
rect 106 -49 107 -48
rect 107 -49 108 -48
rect 108 -49 109 -48
rect 109 -49 110 -48
rect 110 -49 111 -48
rect 111 -49 112 -48
rect 112 -49 113 -48
rect 113 -49 114 -48
rect 114 -49 115 -48
rect 115 -49 116 -48
rect 116 -49 117 -48
rect 117 -49 118 -48
rect 118 -49 119 -48
rect 119 -49 120 -48
rect 120 -49 121 -48
rect 121 -49 122 -48
rect 122 -49 123 -48
rect 123 -49 124 -48
rect 124 -49 125 -48
rect 125 -49 126 -48
rect 126 -49 127 -48
rect 131 -49 132 -48
rect 132 -49 133 -48
rect 133 -49 134 -48
rect 134 -49 135 -48
rect 135 -49 136 -48
rect 136 -49 137 -48
rect 137 -49 138 -48
rect 138 -49 139 -48
rect 139 -49 140 -48
rect 140 -49 141 -48
rect 141 -49 142 -48
rect 142 -49 143 -48
rect 143 -49 144 -48
rect 144 -49 145 -48
rect 145 -49 146 -48
rect 146 -49 147 -48
rect 147 -49 148 -48
rect 148 -49 149 -48
rect 149 -49 150 -48
rect 150 -49 151 -48
rect 151 -49 152 -48
rect 152 -49 153 -48
rect 153 -49 154 -48
rect 154 -49 155 -48
rect 155 -49 156 -48
rect 156 -49 157 -48
rect 157 -49 158 -48
rect 158 -49 159 -48
rect 163 -49 164 -48
rect 164 -49 165 -48
rect 165 -49 166 -48
rect 166 -49 167 -48
rect 167 -49 168 -48
rect 168 -49 169 -48
rect 169 -49 170 -48
rect 170 -49 171 -48
rect 171 -49 172 -48
rect 172 -49 173 -48
rect 173 -49 174 -48
rect 174 -49 175 -48
rect 175 -49 176 -48
rect 176 -49 177 -48
rect 177 -49 178 -48
rect 178 -49 179 -48
rect 179 -49 180 -48
rect 180 -49 181 -48
rect 181 -49 182 -48
rect 182 -49 183 -48
rect 183 -49 184 -48
rect 184 -49 185 -48
rect 185 -49 186 -48
rect 186 -49 187 -48
rect 187 -49 188 -48
rect 188 -49 189 -48
rect 189 -49 190 -48
rect 190 -49 191 -48
rect 191 -49 192 -48
rect 192 -49 193 -48
rect 193 -49 194 -48
rect 194 -49 195 -48
rect 195 -49 196 -48
rect 196 -49 197 -48
rect 197 -49 198 -48
rect 198 -49 199 -48
rect 199 -49 200 -48
rect 200 -49 201 -48
rect 201 -49 202 -48
rect 202 -49 203 -48
rect 203 -49 204 -48
rect 204 -49 205 -48
rect 205 -49 206 -48
rect 206 -49 207 -48
rect 207 -49 208 -48
rect 208 -49 209 -48
rect 209 -49 210 -48
rect 210 -49 211 -48
rect 211 -49 212 -48
rect 212 -49 213 -48
rect 213 -49 214 -48
rect 214 -49 215 -48
rect 215 -49 216 -48
rect 216 -49 217 -48
rect 217 -49 218 -48
rect 218 -49 219 -48
rect 219 -49 220 -48
rect 220 -49 221 -48
rect 221 -49 222 -48
rect 222 -49 223 -48
rect 223 -49 224 -48
rect 224 -49 225 -48
rect 225 -49 226 -48
rect 226 -49 227 -48
rect 227 -49 228 -48
rect 228 -49 229 -48
rect 229 -49 230 -48
rect 230 -49 231 -48
rect 231 -49 232 -48
rect 232 -49 233 -48
rect 233 -49 234 -48
rect 234 -49 235 -48
rect 235 -49 236 -48
rect 236 -49 237 -48
rect 237 -49 238 -48
rect 238 -49 239 -48
rect 239 -49 240 -48
rect 240 -49 241 -48
rect 241 -49 242 -48
rect 242 -49 243 -48
rect 243 -49 244 -48
rect 244 -49 245 -48
rect 245 -49 246 -48
rect 246 -49 247 -48
rect 247 -49 248 -48
rect 248 -49 249 -48
rect 249 -49 250 -48
rect 250 -49 251 -48
rect 251 -49 252 -48
rect 252 -49 253 -48
rect 253 -49 254 -48
rect 254 -49 255 -48
rect 255 -49 256 -48
rect 256 -49 257 -48
rect 257 -49 258 -48
rect 258 -49 259 -48
rect 259 -49 260 -48
rect 260 -49 261 -48
rect 261 -49 262 -48
rect 262 -49 263 -48
rect 263 -49 264 -48
rect 264 -49 265 -48
rect 265 -49 266 -48
rect 266 -49 267 -48
rect 267 -49 268 -48
rect 268 -49 269 -48
rect 269 -49 270 -48
rect 270 -49 271 -48
rect 271 -49 272 -48
rect 272 -49 273 -48
rect 273 -49 274 -48
rect 274 -49 275 -48
rect 275 -49 276 -48
rect 276 -49 277 -48
rect 277 -49 278 -48
rect 278 -49 279 -48
rect 279 -49 280 -48
rect 280 -49 281 -48
rect 281 -49 282 -48
rect 282 -49 283 -48
rect 283 -49 284 -48
rect 284 -49 285 -48
rect 285 -49 286 -48
rect 286 -49 287 -48
rect 287 -49 288 -48
rect 288 -49 289 -48
rect 289 -49 290 -48
rect 290 -49 291 -48
rect 291 -49 292 -48
rect 292 -49 293 -48
rect 293 -49 294 -48
rect 294 -49 295 -48
rect 295 -49 296 -48
rect 296 -49 297 -48
rect 297 -49 298 -48
rect 298 -49 299 -48
rect 299 -49 300 -48
rect 300 -49 301 -48
rect 301 -49 302 -48
rect 302 -49 303 -48
rect 303 -49 304 -48
rect 304 -49 305 -48
rect 305 -49 306 -48
rect 306 -49 307 -48
rect 307 -49 308 -48
rect 308 -49 309 -48
rect 309 -49 310 -48
rect 310 -49 311 -48
rect 311 -49 312 -48
rect 312 -49 313 -48
rect 313 -49 314 -48
rect 314 -49 315 -48
rect 315 -49 316 -48
rect 316 -49 317 -48
rect 317 -49 318 -48
rect 318 -49 319 -48
rect 319 -49 320 -48
rect 320 -49 321 -48
rect 321 -49 322 -48
rect 322 -49 323 -48
rect 323 -49 324 -48
rect 324 -49 325 -48
rect 325 -49 326 -48
rect 326 -49 327 -48
rect 327 -49 328 -48
rect 328 -49 329 -48
rect 329 -49 330 -48
rect 330 -49 331 -48
rect 331 -49 332 -48
rect 332 -49 333 -48
rect 333 -49 334 -48
rect 334 -49 335 -48
rect 335 -49 336 -48
rect 336 -49 337 -48
rect 337 -49 338 -48
rect 338 -49 339 -48
rect 339 -49 340 -48
rect 340 -49 341 -48
rect 341 -49 342 -48
rect 342 -49 343 -48
rect 343 -49 344 -48
rect 344 -49 345 -48
rect 345 -49 346 -48
rect 346 -49 347 -48
rect 347 -49 348 -48
rect 348 -49 349 -48
rect 349 -49 350 -48
rect 350 -49 351 -48
rect 351 -49 352 -48
rect 352 -49 353 -48
rect 353 -49 354 -48
rect 354 -49 355 -48
rect 355 -49 356 -48
rect 356 -49 357 -48
rect 357 -49 358 -48
rect 358 -49 359 -48
rect 359 -49 360 -48
rect 360 -49 361 -48
rect 361 -49 362 -48
rect 362 -49 363 -48
rect 363 -49 364 -48
rect 364 -49 365 -48
rect 365 -49 366 -48
rect 366 -49 367 -48
rect 367 -49 368 -48
rect 368 -49 369 -48
rect 369 -49 370 -48
rect 370 -49 371 -48
rect 371 -49 372 -48
rect 372 -49 373 -48
rect 373 -49 374 -48
rect 374 -49 375 -48
rect 375 -49 376 -48
rect 376 -49 377 -48
rect 377 -49 378 -48
rect 378 -49 379 -48
rect 379 -49 380 -48
rect 380 -49 381 -48
rect 381 -49 382 -48
rect 382 -49 383 -48
rect 383 -49 384 -48
rect 384 -49 385 -48
rect 385 -49 386 -48
rect 386 -49 387 -48
rect 387 -49 388 -48
rect 388 -49 389 -48
rect 389 -49 390 -48
rect 390 -49 391 -48
rect 391 -49 392 -48
rect 392 -49 393 -48
rect 393 -49 394 -48
rect 394 -49 395 -48
rect 395 -49 396 -48
rect 396 -49 397 -48
rect 397 -49 398 -48
rect 398 -49 399 -48
rect 399 -49 400 -48
rect 400 -49 401 -48
rect 401 -49 402 -48
rect 402 -49 403 -48
rect 403 -49 404 -48
rect 404 -49 405 -48
rect 405 -49 406 -48
rect 406 -49 407 -48
rect 407 -49 408 -48
rect 408 -49 409 -48
rect 409 -49 410 -48
rect 410 -49 411 -48
rect 411 -49 412 -48
rect 412 -49 413 -48
rect 413 -49 414 -48
rect 414 -49 415 -48
rect 415 -49 416 -48
rect 416 -49 417 -48
rect 417 -49 418 -48
rect 418 -49 419 -48
rect 419 -49 420 -48
rect 420 -49 421 -48
rect 421 -49 422 -48
rect 422 -49 423 -48
rect 423 -49 424 -48
rect 424 -49 425 -48
rect 425 -49 426 -48
rect 426 -49 427 -48
rect 427 -49 428 -48
rect 428 -49 429 -48
rect 429 -49 430 -48
rect 430 -49 431 -48
rect 431 -49 432 -48
rect 432 -49 433 -48
rect 433 -49 434 -48
rect 434 -49 435 -48
rect 435 -49 436 -48
rect 436 -49 437 -48
rect 437 -49 438 -48
rect 438 -49 439 -48
rect 439 -49 440 -48
rect 440 -49 441 -48
rect 441 -49 442 -48
rect 442 -49 443 -48
rect 443 -49 444 -48
rect 444 -49 445 -48
rect 445 -49 446 -48
rect 446 -49 447 -48
rect 447 -49 448 -48
rect 448 -49 449 -48
rect 449 -49 450 -48
rect 450 -49 451 -48
rect 451 -49 452 -48
rect 452 -49 453 -48
rect 453 -49 454 -48
rect 454 -49 455 -48
rect 455 -49 456 -48
rect 456 -49 457 -48
rect 457 -49 458 -48
rect 458 -49 459 -48
rect 459 -49 460 -48
rect 460 -49 461 -48
rect 461 -49 462 -48
rect 462 -49 463 -48
rect 463 -49 464 -48
rect 464 -49 465 -48
rect 465 -49 466 -48
rect 466 -49 467 -48
rect 467 -49 468 -48
rect 468 -49 469 -48
rect 469 -49 470 -48
rect 470 -49 471 -48
rect 471 -49 472 -48
rect 472 -49 473 -48
rect 473 -49 474 -48
rect 474 -49 475 -48
rect 475 -49 476 -48
rect 476 -49 477 -48
rect 477 -49 478 -48
rect 478 -49 479 -48
rect 479 -49 480 -48
rect 2 -50 3 -49
rect 3 -50 4 -49
rect 4 -50 5 -49
rect 5 -50 6 -49
rect 6 -50 7 -49
rect 7 -50 8 -49
rect 8 -50 9 -49
rect 9 -50 10 -49
rect 10 -50 11 -49
rect 11 -50 12 -49
rect 12 -50 13 -49
rect 13 -50 14 -49
rect 14 -50 15 -49
rect 15 -50 16 -49
rect 16 -50 17 -49
rect 17 -50 18 -49
rect 18 -50 19 -49
rect 19 -50 20 -49
rect 20 -50 21 -49
rect 21 -50 22 -49
rect 22 -50 23 -49
rect 23 -50 24 -49
rect 24 -50 25 -49
rect 25 -50 26 -49
rect 26 -50 27 -49
rect 27 -50 28 -49
rect 28 -50 29 -49
rect 29 -50 30 -49
rect 35 -50 36 -49
rect 36 -50 37 -49
rect 37 -50 38 -49
rect 38 -50 39 -49
rect 39 -50 40 -49
rect 40 -50 41 -49
rect 41 -50 42 -49
rect 42 -50 43 -49
rect 43 -50 44 -49
rect 44 -50 45 -49
rect 45 -50 46 -49
rect 46 -50 47 -49
rect 47 -50 48 -49
rect 48 -50 49 -49
rect 49 -50 50 -49
rect 50 -50 51 -49
rect 51 -50 52 -49
rect 52 -50 53 -49
rect 53 -50 54 -49
rect 54 -50 55 -49
rect 55 -50 56 -49
rect 56 -50 57 -49
rect 57 -50 58 -49
rect 58 -50 59 -49
rect 59 -50 60 -49
rect 60 -50 61 -49
rect 61 -50 62 -49
rect 67 -50 68 -49
rect 68 -50 69 -49
rect 69 -50 70 -49
rect 70 -50 71 -49
rect 71 -50 72 -49
rect 72 -50 73 -49
rect 73 -50 74 -49
rect 74 -50 75 -49
rect 75 -50 76 -49
rect 76 -50 77 -49
rect 77 -50 78 -49
rect 78 -50 79 -49
rect 79 -50 80 -49
rect 80 -50 81 -49
rect 81 -50 82 -49
rect 82 -50 83 -49
rect 83 -50 84 -49
rect 84 -50 85 -49
rect 85 -50 86 -49
rect 86 -50 87 -49
rect 87 -50 88 -49
rect 88 -50 89 -49
rect 89 -50 90 -49
rect 90 -50 91 -49
rect 91 -50 92 -49
rect 92 -50 93 -49
rect 93 -50 94 -49
rect 99 -50 100 -49
rect 100 -50 101 -49
rect 101 -50 102 -49
rect 102 -50 103 -49
rect 103 -50 104 -49
rect 104 -50 105 -49
rect 105 -50 106 -49
rect 106 -50 107 -49
rect 107 -50 108 -49
rect 108 -50 109 -49
rect 109 -50 110 -49
rect 110 -50 111 -49
rect 111 -50 112 -49
rect 112 -50 113 -49
rect 113 -50 114 -49
rect 114 -50 115 -49
rect 115 -50 116 -49
rect 116 -50 117 -49
rect 117 -50 118 -49
rect 118 -50 119 -49
rect 119 -50 120 -49
rect 120 -50 121 -49
rect 121 -50 122 -49
rect 122 -50 123 -49
rect 123 -50 124 -49
rect 124 -50 125 -49
rect 125 -50 126 -49
rect 131 -50 132 -49
rect 132 -50 133 -49
rect 133 -50 134 -49
rect 134 -50 135 -49
rect 135 -50 136 -49
rect 136 -50 137 -49
rect 137 -50 138 -49
rect 138 -50 139 -49
rect 139 -50 140 -49
rect 140 -50 141 -49
rect 141 -50 142 -49
rect 142 -50 143 -49
rect 143 -50 144 -49
rect 144 -50 145 -49
rect 145 -50 146 -49
rect 146 -50 147 -49
rect 147 -50 148 -49
rect 148 -50 149 -49
rect 149 -50 150 -49
rect 150 -50 151 -49
rect 151 -50 152 -49
rect 152 -50 153 -49
rect 153 -50 154 -49
rect 154 -50 155 -49
rect 155 -50 156 -49
rect 156 -50 157 -49
rect 157 -50 158 -49
rect 163 -50 164 -49
rect 164 -50 165 -49
rect 165 -50 166 -49
rect 166 -50 167 -49
rect 167 -50 168 -49
rect 168 -50 169 -49
rect 169 -50 170 -49
rect 170 -50 171 -49
rect 171 -50 172 -49
rect 172 -50 173 -49
rect 173 -50 174 -49
rect 174 -50 175 -49
rect 175 -50 176 -49
rect 176 -50 177 -49
rect 177 -50 178 -49
rect 178 -50 179 -49
rect 179 -50 180 -49
rect 180 -50 181 -49
rect 181 -50 182 -49
rect 182 -50 183 -49
rect 183 -50 184 -49
rect 184 -50 185 -49
rect 185 -50 186 -49
rect 186 -50 187 -49
rect 187 -50 188 -49
rect 188 -50 189 -49
rect 189 -50 190 -49
rect 190 -50 191 -49
rect 191 -50 192 -49
rect 192 -50 193 -49
rect 193 -50 194 -49
rect 194 -50 195 -49
rect 195 -50 196 -49
rect 196 -50 197 -49
rect 197 -50 198 -49
rect 198 -50 199 -49
rect 199 -50 200 -49
rect 200 -50 201 -49
rect 201 -50 202 -49
rect 202 -50 203 -49
rect 203 -50 204 -49
rect 204 -50 205 -49
rect 205 -50 206 -49
rect 206 -50 207 -49
rect 207 -50 208 -49
rect 208 -50 209 -49
rect 209 -50 210 -49
rect 210 -50 211 -49
rect 211 -50 212 -49
rect 212 -50 213 -49
rect 213 -50 214 -49
rect 214 -50 215 -49
rect 215 -50 216 -49
rect 216 -50 217 -49
rect 217 -50 218 -49
rect 218 -50 219 -49
rect 219 -50 220 -49
rect 220 -50 221 -49
rect 221 -50 222 -49
rect 222 -50 223 -49
rect 223 -50 224 -49
rect 224 -50 225 -49
rect 225 -50 226 -49
rect 226 -50 227 -49
rect 227 -50 228 -49
rect 228 -50 229 -49
rect 229 -50 230 -49
rect 230 -50 231 -49
rect 231 -50 232 -49
rect 232 -50 233 -49
rect 233 -50 234 -49
rect 234 -50 235 -49
rect 235 -50 236 -49
rect 236 -50 237 -49
rect 237 -50 238 -49
rect 238 -50 239 -49
rect 239 -50 240 -49
rect 240 -50 241 -49
rect 241 -50 242 -49
rect 242 -50 243 -49
rect 243 -50 244 -49
rect 244 -50 245 -49
rect 245 -50 246 -49
rect 246 -50 247 -49
rect 247 -50 248 -49
rect 248 -50 249 -49
rect 249 -50 250 -49
rect 250 -50 251 -49
rect 251 -50 252 -49
rect 252 -50 253 -49
rect 253 -50 254 -49
rect 254 -50 255 -49
rect 255 -50 256 -49
rect 256 -50 257 -49
rect 257 -50 258 -49
rect 258 -50 259 -49
rect 259 -50 260 -49
rect 260 -50 261 -49
rect 261 -50 262 -49
rect 262 -50 263 -49
rect 263 -50 264 -49
rect 264 -50 265 -49
rect 265 -50 266 -49
rect 266 -50 267 -49
rect 267 -50 268 -49
rect 268 -50 269 -49
rect 269 -50 270 -49
rect 270 -50 271 -49
rect 271 -50 272 -49
rect 272 -50 273 -49
rect 273 -50 274 -49
rect 274 -50 275 -49
rect 275 -50 276 -49
rect 276 -50 277 -49
rect 277 -50 278 -49
rect 278 -50 279 -49
rect 279 -50 280 -49
rect 280 -50 281 -49
rect 281 -50 282 -49
rect 282 -50 283 -49
rect 283 -50 284 -49
rect 284 -50 285 -49
rect 285 -50 286 -49
rect 286 -50 287 -49
rect 287 -50 288 -49
rect 288 -50 289 -49
rect 289 -50 290 -49
rect 290 -50 291 -49
rect 291 -50 292 -49
rect 292 -50 293 -49
rect 293 -50 294 -49
rect 294 -50 295 -49
rect 295 -50 296 -49
rect 296 -50 297 -49
rect 297 -50 298 -49
rect 298 -50 299 -49
rect 299 -50 300 -49
rect 300 -50 301 -49
rect 301 -50 302 -49
rect 302 -50 303 -49
rect 303 -50 304 -49
rect 304 -50 305 -49
rect 305 -50 306 -49
rect 306 -50 307 -49
rect 307 -50 308 -49
rect 308 -50 309 -49
rect 309 -50 310 -49
rect 310 -50 311 -49
rect 311 -50 312 -49
rect 312 -50 313 -49
rect 313 -50 314 -49
rect 314 -50 315 -49
rect 315 -50 316 -49
rect 316 -50 317 -49
rect 317 -50 318 -49
rect 318 -50 319 -49
rect 319 -50 320 -49
rect 320 -50 321 -49
rect 321 -50 322 -49
rect 322 -50 323 -49
rect 323 -50 324 -49
rect 324 -50 325 -49
rect 325 -50 326 -49
rect 326 -50 327 -49
rect 327 -50 328 -49
rect 328 -50 329 -49
rect 329 -50 330 -49
rect 330 -50 331 -49
rect 331 -50 332 -49
rect 332 -50 333 -49
rect 333 -50 334 -49
rect 334 -50 335 -49
rect 335 -50 336 -49
rect 336 -50 337 -49
rect 337 -50 338 -49
rect 338 -50 339 -49
rect 339 -50 340 -49
rect 340 -50 341 -49
rect 341 -50 342 -49
rect 342 -50 343 -49
rect 343 -50 344 -49
rect 344 -50 345 -49
rect 345 -50 346 -49
rect 346 -50 347 -49
rect 347 -50 348 -49
rect 348 -50 349 -49
rect 349 -50 350 -49
rect 350 -50 351 -49
rect 351 -50 352 -49
rect 352 -50 353 -49
rect 353 -50 354 -49
rect 354 -50 355 -49
rect 355 -50 356 -49
rect 356 -50 357 -49
rect 357 -50 358 -49
rect 358 -50 359 -49
rect 359 -50 360 -49
rect 360 -50 361 -49
rect 361 -50 362 -49
rect 362 -50 363 -49
rect 363 -50 364 -49
rect 364 -50 365 -49
rect 365 -50 366 -49
rect 366 -50 367 -49
rect 367 -50 368 -49
rect 368 -50 369 -49
rect 369 -50 370 -49
rect 370 -50 371 -49
rect 371 -50 372 -49
rect 372 -50 373 -49
rect 373 -50 374 -49
rect 374 -50 375 -49
rect 375 -50 376 -49
rect 376 -50 377 -49
rect 377 -50 378 -49
rect 378 -50 379 -49
rect 379 -50 380 -49
rect 380 -50 381 -49
rect 381 -50 382 -49
rect 382 -50 383 -49
rect 383 -50 384 -49
rect 384 -50 385 -49
rect 385 -50 386 -49
rect 386 -50 387 -49
rect 387 -50 388 -49
rect 388 -50 389 -49
rect 389 -50 390 -49
rect 390 -50 391 -49
rect 391 -50 392 -49
rect 392 -50 393 -49
rect 393 -50 394 -49
rect 394 -50 395 -49
rect 395 -50 396 -49
rect 396 -50 397 -49
rect 397 -50 398 -49
rect 398 -50 399 -49
rect 399 -50 400 -49
rect 400 -50 401 -49
rect 401 -50 402 -49
rect 402 -50 403 -49
rect 403 -50 404 -49
rect 404 -50 405 -49
rect 405 -50 406 -49
rect 406 -50 407 -49
rect 407 -50 408 -49
rect 408 -50 409 -49
rect 409 -50 410 -49
rect 410 -50 411 -49
rect 411 -50 412 -49
rect 412 -50 413 -49
rect 413 -50 414 -49
rect 414 -50 415 -49
rect 415 -50 416 -49
rect 416 -50 417 -49
rect 417 -50 418 -49
rect 418 -50 419 -49
rect 419 -50 420 -49
rect 420 -50 421 -49
rect 421 -50 422 -49
rect 422 -50 423 -49
rect 423 -50 424 -49
rect 424 -50 425 -49
rect 425 -50 426 -49
rect 426 -50 427 -49
rect 427 -50 428 -49
rect 428 -50 429 -49
rect 429 -50 430 -49
rect 430 -50 431 -49
rect 431 -50 432 -49
rect 432 -50 433 -49
rect 433 -50 434 -49
rect 434 -50 435 -49
rect 435 -50 436 -49
rect 436 -50 437 -49
rect 437 -50 438 -49
rect 438 -50 439 -49
rect 439 -50 440 -49
rect 440 -50 441 -49
rect 441 -50 442 -49
rect 442 -50 443 -49
rect 443 -50 444 -49
rect 444 -50 445 -49
rect 445 -50 446 -49
rect 446 -50 447 -49
rect 447 -50 448 -49
rect 448 -50 449 -49
rect 449 -50 450 -49
rect 450 -50 451 -49
rect 451 -50 452 -49
rect 452 -50 453 -49
rect 453 -50 454 -49
rect 454 -50 455 -49
rect 455 -50 456 -49
rect 456 -50 457 -49
rect 457 -50 458 -49
rect 458 -50 459 -49
rect 459 -50 460 -49
rect 460 -50 461 -49
rect 461 -50 462 -49
rect 462 -50 463 -49
rect 463 -50 464 -49
rect 464 -50 465 -49
rect 465 -50 466 -49
rect 466 -50 467 -49
rect 467 -50 468 -49
rect 468 -50 469 -49
rect 469 -50 470 -49
rect 470 -50 471 -49
rect 471 -50 472 -49
rect 472 -50 473 -49
rect 473 -50 474 -49
rect 474 -50 475 -49
rect 475 -50 476 -49
rect 476 -50 477 -49
rect 477 -50 478 -49
rect 478 -50 479 -49
rect 479 -50 480 -49
rect 2 -51 3 -50
rect 3 -51 4 -50
rect 4 -51 5 -50
rect 5 -51 6 -50
rect 6 -51 7 -50
rect 7 -51 8 -50
rect 8 -51 9 -50
rect 9 -51 10 -50
rect 10 -51 11 -50
rect 11 -51 12 -50
rect 12 -51 13 -50
rect 13 -51 14 -50
rect 14 -51 15 -50
rect 15 -51 16 -50
rect 16 -51 17 -50
rect 17 -51 18 -50
rect 18 -51 19 -50
rect 19 -51 20 -50
rect 20 -51 21 -50
rect 21 -51 22 -50
rect 22 -51 23 -50
rect 23 -51 24 -50
rect 24 -51 25 -50
rect 41 -51 42 -50
rect 42 -51 43 -50
rect 43 -51 44 -50
rect 44 -51 45 -50
rect 45 -51 46 -50
rect 46 -51 47 -50
rect 47 -51 48 -50
rect 48 -51 49 -50
rect 49 -51 50 -50
rect 50 -51 51 -50
rect 51 -51 52 -50
rect 52 -51 53 -50
rect 53 -51 54 -50
rect 54 -51 55 -50
rect 55 -51 56 -50
rect 56 -51 57 -50
rect 73 -51 74 -50
rect 74 -51 75 -50
rect 75 -51 76 -50
rect 76 -51 77 -50
rect 77 -51 78 -50
rect 78 -51 79 -50
rect 79 -51 80 -50
rect 80 -51 81 -50
rect 81 -51 82 -50
rect 82 -51 83 -50
rect 83 -51 84 -50
rect 84 -51 85 -50
rect 85 -51 86 -50
rect 86 -51 87 -50
rect 87 -51 88 -50
rect 88 -51 89 -50
rect 105 -51 106 -50
rect 106 -51 107 -50
rect 107 -51 108 -50
rect 108 -51 109 -50
rect 109 -51 110 -50
rect 110 -51 111 -50
rect 111 -51 112 -50
rect 112 -51 113 -50
rect 113 -51 114 -50
rect 114 -51 115 -50
rect 115 -51 116 -50
rect 116 -51 117 -50
rect 117 -51 118 -50
rect 118 -51 119 -50
rect 119 -51 120 -50
rect 120 -51 121 -50
rect 137 -51 138 -50
rect 138 -51 139 -50
rect 139 -51 140 -50
rect 140 -51 141 -50
rect 141 -51 142 -50
rect 142 -51 143 -50
rect 143 -51 144 -50
rect 144 -51 145 -50
rect 145 -51 146 -50
rect 146 -51 147 -50
rect 147 -51 148 -50
rect 148 -51 149 -50
rect 149 -51 150 -50
rect 150 -51 151 -50
rect 151 -51 152 -50
rect 152 -51 153 -50
rect 169 -51 170 -50
rect 170 -51 171 -50
rect 171 -51 172 -50
rect 172 -51 173 -50
rect 173 -51 174 -50
rect 174 -51 175 -50
rect 175 -51 176 -50
rect 176 -51 177 -50
rect 177 -51 178 -50
rect 178 -51 179 -50
rect 179 -51 180 -50
rect 180 -51 181 -50
rect 181 -51 182 -50
rect 182 -51 183 -50
rect 183 -51 184 -50
rect 184 -51 185 -50
rect 185 -51 186 -50
rect 186 -51 187 -50
rect 187 -51 188 -50
rect 188 -51 189 -50
rect 189 -51 190 -50
rect 190 -51 191 -50
rect 191 -51 192 -50
rect 192 -51 193 -50
rect 193 -51 194 -50
rect 194 -51 195 -50
rect 195 -51 196 -50
rect 196 -51 197 -50
rect 197 -51 198 -50
rect 198 -51 199 -50
rect 199 -51 200 -50
rect 200 -51 201 -50
rect 201 -51 202 -50
rect 202 -51 203 -50
rect 203 -51 204 -50
rect 204 -51 205 -50
rect 205 -51 206 -50
rect 206 -51 207 -50
rect 207 -51 208 -50
rect 208 -51 209 -50
rect 209 -51 210 -50
rect 210 -51 211 -50
rect 211 -51 212 -50
rect 212 -51 213 -50
rect 213 -51 214 -50
rect 214 -51 215 -50
rect 215 -51 216 -50
rect 216 -51 217 -50
rect 217 -51 218 -50
rect 218 -51 219 -50
rect 219 -51 220 -50
rect 220 -51 221 -50
rect 221 -51 222 -50
rect 222 -51 223 -50
rect 223 -51 224 -50
rect 224 -51 225 -50
rect 225 -51 226 -50
rect 226 -51 227 -50
rect 227 -51 228 -50
rect 228 -51 229 -50
rect 229 -51 230 -50
rect 230 -51 231 -50
rect 231 -51 232 -50
rect 232 -51 233 -50
rect 233 -51 234 -50
rect 234 -51 235 -50
rect 235 -51 236 -50
rect 236 -51 237 -50
rect 237 -51 238 -50
rect 238 -51 239 -50
rect 239 -51 240 -50
rect 240 -51 241 -50
rect 241 -51 242 -50
rect 242 -51 243 -50
rect 243 -51 244 -50
rect 244 -51 245 -50
rect 245 -51 246 -50
rect 246 -51 247 -50
rect 247 -51 248 -50
rect 248 -51 249 -50
rect 249 -51 250 -50
rect 250 -51 251 -50
rect 251 -51 252 -50
rect 252 -51 253 -50
rect 253 -51 254 -50
rect 254 -51 255 -50
rect 255 -51 256 -50
rect 256 -51 257 -50
rect 257 -51 258 -50
rect 258 -51 259 -50
rect 259 -51 260 -50
rect 260 -51 261 -50
rect 261 -51 262 -50
rect 262 -51 263 -50
rect 263 -51 264 -50
rect 264 -51 265 -50
rect 265 -51 266 -50
rect 266 -51 267 -50
rect 267 -51 268 -50
rect 268 -51 269 -50
rect 269 -51 270 -50
rect 270 -51 271 -50
rect 271 -51 272 -50
rect 272 -51 273 -50
rect 273 -51 274 -50
rect 274 -51 275 -50
rect 275 -51 276 -50
rect 276 -51 277 -50
rect 277 -51 278 -50
rect 278 -51 279 -50
rect 279 -51 280 -50
rect 280 -51 281 -50
rect 281 -51 282 -50
rect 282 -51 283 -50
rect 283 -51 284 -50
rect 284 -51 285 -50
rect 285 -51 286 -50
rect 286 -51 287 -50
rect 287 -51 288 -50
rect 288 -51 289 -50
rect 289 -51 290 -50
rect 290 -51 291 -50
rect 291 -51 292 -50
rect 292 -51 293 -50
rect 293 -51 294 -50
rect 294 -51 295 -50
rect 295 -51 296 -50
rect 296 -51 297 -50
rect 297 -51 298 -50
rect 298 -51 299 -50
rect 299 -51 300 -50
rect 300 -51 301 -50
rect 301 -51 302 -50
rect 302 -51 303 -50
rect 303 -51 304 -50
rect 304 -51 305 -50
rect 305 -51 306 -50
rect 306 -51 307 -50
rect 307 -51 308 -50
rect 308 -51 309 -50
rect 309 -51 310 -50
rect 310 -51 311 -50
rect 311 -51 312 -50
rect 312 -51 313 -50
rect 313 -51 314 -50
rect 314 -51 315 -50
rect 315 -51 316 -50
rect 316 -51 317 -50
rect 317 -51 318 -50
rect 318 -51 319 -50
rect 319 -51 320 -50
rect 320 -51 321 -50
rect 321 -51 322 -50
rect 322 -51 323 -50
rect 323 -51 324 -50
rect 324 -51 325 -50
rect 325 -51 326 -50
rect 326 -51 327 -50
rect 327 -51 328 -50
rect 328 -51 329 -50
rect 329 -51 330 -50
rect 330 -51 331 -50
rect 331 -51 332 -50
rect 332 -51 333 -50
rect 333 -51 334 -50
rect 334 -51 335 -50
rect 335 -51 336 -50
rect 336 -51 337 -50
rect 337 -51 338 -50
rect 338 -51 339 -50
rect 339 -51 340 -50
rect 340 -51 341 -50
rect 341 -51 342 -50
rect 342 -51 343 -50
rect 343 -51 344 -50
rect 344 -51 345 -50
rect 345 -51 346 -50
rect 346 -51 347 -50
rect 347 -51 348 -50
rect 348 -51 349 -50
rect 349 -51 350 -50
rect 350 -51 351 -50
rect 351 -51 352 -50
rect 352 -51 353 -50
rect 353 -51 354 -50
rect 354 -51 355 -50
rect 355 -51 356 -50
rect 356 -51 357 -50
rect 357 -51 358 -50
rect 358 -51 359 -50
rect 359 -51 360 -50
rect 360 -51 361 -50
rect 361 -51 362 -50
rect 362 -51 363 -50
rect 363 -51 364 -50
rect 364 -51 365 -50
rect 365 -51 366 -50
rect 366 -51 367 -50
rect 367 -51 368 -50
rect 368 -51 369 -50
rect 369 -51 370 -50
rect 370 -51 371 -50
rect 371 -51 372 -50
rect 372 -51 373 -50
rect 373 -51 374 -50
rect 374 -51 375 -50
rect 375 -51 376 -50
rect 376 -51 377 -50
rect 377 -51 378 -50
rect 378 -51 379 -50
rect 379 -51 380 -50
rect 380 -51 381 -50
rect 381 -51 382 -50
rect 382 -51 383 -50
rect 383 -51 384 -50
rect 384 -51 385 -50
rect 385 -51 386 -50
rect 386 -51 387 -50
rect 387 -51 388 -50
rect 388 -51 389 -50
rect 389 -51 390 -50
rect 390 -51 391 -50
rect 391 -51 392 -50
rect 392 -51 393 -50
rect 393 -51 394 -50
rect 394 -51 395 -50
rect 395 -51 396 -50
rect 396 -51 397 -50
rect 397 -51 398 -50
rect 398 -51 399 -50
rect 399 -51 400 -50
rect 400 -51 401 -50
rect 401 -51 402 -50
rect 402 -51 403 -50
rect 403 -51 404 -50
rect 404 -51 405 -50
rect 405 -51 406 -50
rect 406 -51 407 -50
rect 407 -51 408 -50
rect 408 -51 409 -50
rect 409 -51 410 -50
rect 410 -51 411 -50
rect 411 -51 412 -50
rect 412 -51 413 -50
rect 413 -51 414 -50
rect 414 -51 415 -50
rect 415 -51 416 -50
rect 416 -51 417 -50
rect 417 -51 418 -50
rect 418 -51 419 -50
rect 419 -51 420 -50
rect 420 -51 421 -50
rect 421 -51 422 -50
rect 422 -51 423 -50
rect 423 -51 424 -50
rect 424 -51 425 -50
rect 425 -51 426 -50
rect 426 -51 427 -50
rect 427 -51 428 -50
rect 428 -51 429 -50
rect 429 -51 430 -50
rect 430 -51 431 -50
rect 431 -51 432 -50
rect 432 -51 433 -50
rect 433 -51 434 -50
rect 434 -51 435 -50
rect 435 -51 436 -50
rect 436 -51 437 -50
rect 437 -51 438 -50
rect 438 -51 439 -50
rect 439 -51 440 -50
rect 440 -51 441 -50
rect 441 -51 442 -50
rect 442 -51 443 -50
rect 443 -51 444 -50
rect 444 -51 445 -50
rect 445 -51 446 -50
rect 446 -51 447 -50
rect 447 -51 448 -50
rect 448 -51 449 -50
rect 449 -51 450 -50
rect 450 -51 451 -50
rect 451 -51 452 -50
rect 452 -51 453 -50
rect 453 -51 454 -50
rect 454 -51 455 -50
rect 455 -51 456 -50
rect 456 -51 457 -50
rect 457 -51 458 -50
rect 458 -51 459 -50
rect 459 -51 460 -50
rect 460 -51 461 -50
rect 461 -51 462 -50
rect 462 -51 463 -50
rect 463 -51 464 -50
rect 464 -51 465 -50
rect 465 -51 466 -50
rect 466 -51 467 -50
rect 467 -51 468 -50
rect 468 -51 469 -50
rect 469 -51 470 -50
rect 470 -51 471 -50
rect 471 -51 472 -50
rect 472 -51 473 -50
rect 473 -51 474 -50
rect 474 -51 475 -50
rect 475 -51 476 -50
rect 476 -51 477 -50
rect 477 -51 478 -50
rect 478 -51 479 -50
rect 479 -51 480 -50
rect 2 -52 3 -51
rect 3 -52 4 -51
rect 4 -52 5 -51
rect 5 -52 6 -51
rect 6 -52 7 -51
rect 7 -52 8 -51
rect 8 -52 9 -51
rect 9 -52 10 -51
rect 10 -52 11 -51
rect 11 -52 12 -51
rect 12 -52 13 -51
rect 13 -52 14 -51
rect 14 -52 15 -51
rect 15 -52 16 -51
rect 16 -52 17 -51
rect 17 -52 18 -51
rect 18 -52 19 -51
rect 19 -52 20 -51
rect 20 -52 21 -51
rect 21 -52 22 -51
rect 22 -52 23 -51
rect 23 -52 24 -51
rect 24 -52 25 -51
rect 41 -52 42 -51
rect 42 -52 43 -51
rect 43 -52 44 -51
rect 44 -52 45 -51
rect 45 -52 46 -51
rect 46 -52 47 -51
rect 47 -52 48 -51
rect 48 -52 49 -51
rect 49 -52 50 -51
rect 50 -52 51 -51
rect 51 -52 52 -51
rect 52 -52 53 -51
rect 53 -52 54 -51
rect 54 -52 55 -51
rect 55 -52 56 -51
rect 56 -52 57 -51
rect 73 -52 74 -51
rect 74 -52 75 -51
rect 75 -52 76 -51
rect 76 -52 77 -51
rect 77 -52 78 -51
rect 78 -52 79 -51
rect 79 -52 80 -51
rect 80 -52 81 -51
rect 81 -52 82 -51
rect 82 -52 83 -51
rect 83 -52 84 -51
rect 84 -52 85 -51
rect 85 -52 86 -51
rect 86 -52 87 -51
rect 87 -52 88 -51
rect 88 -52 89 -51
rect 105 -52 106 -51
rect 106 -52 107 -51
rect 107 -52 108 -51
rect 108 -52 109 -51
rect 109 -52 110 -51
rect 110 -52 111 -51
rect 111 -52 112 -51
rect 112 -52 113 -51
rect 113 -52 114 -51
rect 114 -52 115 -51
rect 115 -52 116 -51
rect 116 -52 117 -51
rect 117 -52 118 -51
rect 118 -52 119 -51
rect 119 -52 120 -51
rect 120 -52 121 -51
rect 137 -52 138 -51
rect 138 -52 139 -51
rect 139 -52 140 -51
rect 140 -52 141 -51
rect 141 -52 142 -51
rect 142 -52 143 -51
rect 143 -52 144 -51
rect 144 -52 145 -51
rect 145 -52 146 -51
rect 146 -52 147 -51
rect 147 -52 148 -51
rect 148 -52 149 -51
rect 149 -52 150 -51
rect 150 -52 151 -51
rect 151 -52 152 -51
rect 152 -52 153 -51
rect 169 -52 170 -51
rect 170 -52 171 -51
rect 171 -52 172 -51
rect 172 -52 173 -51
rect 173 -52 174 -51
rect 174 -52 175 -51
rect 175 -52 176 -51
rect 176 -52 177 -51
rect 177 -52 178 -51
rect 178 -52 179 -51
rect 179 -52 180 -51
rect 180 -52 181 -51
rect 181 -52 182 -51
rect 182 -52 183 -51
rect 183 -52 184 -51
rect 184 -52 185 -51
rect 185 -52 186 -51
rect 186 -52 187 -51
rect 187 -52 188 -51
rect 188 -52 189 -51
rect 189 -52 190 -51
rect 190 -52 191 -51
rect 191 -52 192 -51
rect 192 -52 193 -51
rect 193 -52 194 -51
rect 194 -52 195 -51
rect 195 -52 196 -51
rect 196 -52 197 -51
rect 197 -52 198 -51
rect 198 -52 199 -51
rect 199 -52 200 -51
rect 200 -52 201 -51
rect 201 -52 202 -51
rect 202 -52 203 -51
rect 203 -52 204 -51
rect 204 -52 205 -51
rect 205 -52 206 -51
rect 206 -52 207 -51
rect 207 -52 208 -51
rect 208 -52 209 -51
rect 209 -52 210 -51
rect 210 -52 211 -51
rect 211 -52 212 -51
rect 212 -52 213 -51
rect 213 -52 214 -51
rect 214 -52 215 -51
rect 215 -52 216 -51
rect 216 -52 217 -51
rect 217 -52 218 -51
rect 218 -52 219 -51
rect 219 -52 220 -51
rect 220 -52 221 -51
rect 221 -52 222 -51
rect 222 -52 223 -51
rect 223 -52 224 -51
rect 224 -52 225 -51
rect 225 -52 226 -51
rect 226 -52 227 -51
rect 227 -52 228 -51
rect 228 -52 229 -51
rect 229 -52 230 -51
rect 230 -52 231 -51
rect 231 -52 232 -51
rect 232 -52 233 -51
rect 233 -52 234 -51
rect 234 -52 235 -51
rect 235 -52 236 -51
rect 236 -52 237 -51
rect 237 -52 238 -51
rect 238 -52 239 -51
rect 239 -52 240 -51
rect 240 -52 241 -51
rect 241 -52 242 -51
rect 242 -52 243 -51
rect 243 -52 244 -51
rect 244 -52 245 -51
rect 245 -52 246 -51
rect 246 -52 247 -51
rect 247 -52 248 -51
rect 248 -52 249 -51
rect 249 -52 250 -51
rect 250 -52 251 -51
rect 251 -52 252 -51
rect 252 -52 253 -51
rect 253 -52 254 -51
rect 254 -52 255 -51
rect 255 -52 256 -51
rect 256 -52 257 -51
rect 257 -52 258 -51
rect 258 -52 259 -51
rect 259 -52 260 -51
rect 260 -52 261 -51
rect 261 -52 262 -51
rect 262 -52 263 -51
rect 263 -52 264 -51
rect 264 -52 265 -51
rect 265 -52 266 -51
rect 266 -52 267 -51
rect 267 -52 268 -51
rect 268 -52 269 -51
rect 269 -52 270 -51
rect 270 -52 271 -51
rect 271 -52 272 -51
rect 272 -52 273 -51
rect 273 -52 274 -51
rect 274 -52 275 -51
rect 275 -52 276 -51
rect 276 -52 277 -51
rect 277 -52 278 -51
rect 278 -52 279 -51
rect 279 -52 280 -51
rect 280 -52 281 -51
rect 281 -52 282 -51
rect 282 -52 283 -51
rect 283 -52 284 -51
rect 284 -52 285 -51
rect 285 -52 286 -51
rect 286 -52 287 -51
rect 287 -52 288 -51
rect 288 -52 289 -51
rect 289 -52 290 -51
rect 290 -52 291 -51
rect 291 -52 292 -51
rect 292 -52 293 -51
rect 293 -52 294 -51
rect 294 -52 295 -51
rect 295 -52 296 -51
rect 296 -52 297 -51
rect 297 -52 298 -51
rect 298 -52 299 -51
rect 299 -52 300 -51
rect 300 -52 301 -51
rect 301 -52 302 -51
rect 302 -52 303 -51
rect 303 -52 304 -51
rect 304 -52 305 -51
rect 305 -52 306 -51
rect 306 -52 307 -51
rect 307 -52 308 -51
rect 308 -52 309 -51
rect 309 -52 310 -51
rect 310 -52 311 -51
rect 311 -52 312 -51
rect 312 -52 313 -51
rect 313 -52 314 -51
rect 314 -52 315 -51
rect 315 -52 316 -51
rect 316 -52 317 -51
rect 317 -52 318 -51
rect 318 -52 319 -51
rect 319 -52 320 -51
rect 320 -52 321 -51
rect 321 -52 322 -51
rect 322 -52 323 -51
rect 323 -52 324 -51
rect 324 -52 325 -51
rect 325 -52 326 -51
rect 326 -52 327 -51
rect 327 -52 328 -51
rect 328 -52 329 -51
rect 329 -52 330 -51
rect 330 -52 331 -51
rect 331 -52 332 -51
rect 332 -52 333 -51
rect 333 -52 334 -51
rect 334 -52 335 -51
rect 335 -52 336 -51
rect 336 -52 337 -51
rect 337 -52 338 -51
rect 338 -52 339 -51
rect 339 -52 340 -51
rect 340 -52 341 -51
rect 341 -52 342 -51
rect 342 -52 343 -51
rect 343 -52 344 -51
rect 344 -52 345 -51
rect 345 -52 346 -51
rect 346 -52 347 -51
rect 347 -52 348 -51
rect 348 -52 349 -51
rect 349 -52 350 -51
rect 350 -52 351 -51
rect 351 -52 352 -51
rect 352 -52 353 -51
rect 353 -52 354 -51
rect 354 -52 355 -51
rect 355 -52 356 -51
rect 356 -52 357 -51
rect 357 -52 358 -51
rect 358 -52 359 -51
rect 359 -52 360 -51
rect 360 -52 361 -51
rect 361 -52 362 -51
rect 362 -52 363 -51
rect 363 -52 364 -51
rect 364 -52 365 -51
rect 365 -52 366 -51
rect 366 -52 367 -51
rect 367 -52 368 -51
rect 368 -52 369 -51
rect 369 -52 370 -51
rect 370 -52 371 -51
rect 371 -52 372 -51
rect 372 -52 373 -51
rect 373 -52 374 -51
rect 374 -52 375 -51
rect 375 -52 376 -51
rect 376 -52 377 -51
rect 377 -52 378 -51
rect 378 -52 379 -51
rect 379 -52 380 -51
rect 380 -52 381 -51
rect 381 -52 382 -51
rect 382 -52 383 -51
rect 383 -52 384 -51
rect 384 -52 385 -51
rect 385 -52 386 -51
rect 386 -52 387 -51
rect 387 -52 388 -51
rect 388 -52 389 -51
rect 389 -52 390 -51
rect 390 -52 391 -51
rect 391 -52 392 -51
rect 392 -52 393 -51
rect 393 -52 394 -51
rect 394 -52 395 -51
rect 395 -52 396 -51
rect 396 -52 397 -51
rect 397 -52 398 -51
rect 398 -52 399 -51
rect 399 -52 400 -51
rect 400 -52 401 -51
rect 401 -52 402 -51
rect 402 -52 403 -51
rect 403 -52 404 -51
rect 404 -52 405 -51
rect 405 -52 406 -51
rect 406 -52 407 -51
rect 407 -52 408 -51
rect 408 -52 409 -51
rect 409 -52 410 -51
rect 410 -52 411 -51
rect 411 -52 412 -51
rect 412 -52 413 -51
rect 413 -52 414 -51
rect 414 -52 415 -51
rect 415 -52 416 -51
rect 416 -52 417 -51
rect 417 -52 418 -51
rect 418 -52 419 -51
rect 419 -52 420 -51
rect 420 -52 421 -51
rect 421 -52 422 -51
rect 422 -52 423 -51
rect 423 -52 424 -51
rect 424 -52 425 -51
rect 425 -52 426 -51
rect 426 -52 427 -51
rect 427 -52 428 -51
rect 428 -52 429 -51
rect 429 -52 430 -51
rect 430 -52 431 -51
rect 431 -52 432 -51
rect 432 -52 433 -51
rect 433 -52 434 -51
rect 434 -52 435 -51
rect 435 -52 436 -51
rect 436 -52 437 -51
rect 437 -52 438 -51
rect 438 -52 439 -51
rect 439 -52 440 -51
rect 440 -52 441 -51
rect 441 -52 442 -51
rect 442 -52 443 -51
rect 443 -52 444 -51
rect 444 -52 445 -51
rect 445 -52 446 -51
rect 446 -52 447 -51
rect 447 -52 448 -51
rect 448 -52 449 -51
rect 449 -52 450 -51
rect 450 -52 451 -51
rect 451 -52 452 -51
rect 452 -52 453 -51
rect 453 -52 454 -51
rect 454 -52 455 -51
rect 455 -52 456 -51
rect 456 -52 457 -51
rect 457 -52 458 -51
rect 458 -52 459 -51
rect 459 -52 460 -51
rect 460 -52 461 -51
rect 461 -52 462 -51
rect 462 -52 463 -51
rect 463 -52 464 -51
rect 464 -52 465 -51
rect 465 -52 466 -51
rect 466 -52 467 -51
rect 467 -52 468 -51
rect 468 -52 469 -51
rect 469 -52 470 -51
rect 470 -52 471 -51
rect 471 -52 472 -51
rect 472 -52 473 -51
rect 473 -52 474 -51
rect 474 -52 475 -51
rect 475 -52 476 -51
rect 476 -52 477 -51
rect 477 -52 478 -51
rect 478 -52 479 -51
rect 479 -52 480 -51
rect 2 -53 3 -52
rect 3 -53 4 -52
rect 4 -53 5 -52
rect 5 -53 6 -52
rect 6 -53 7 -52
rect 7 -53 8 -52
rect 8 -53 9 -52
rect 9 -53 10 -52
rect 10 -53 11 -52
rect 11 -53 12 -52
rect 12 -53 13 -52
rect 13 -53 14 -52
rect 14 -53 15 -52
rect 15 -53 16 -52
rect 16 -53 17 -52
rect 17 -53 18 -52
rect 18 -53 19 -52
rect 19 -53 20 -52
rect 20 -53 21 -52
rect 21 -53 22 -52
rect 22 -53 23 -52
rect 23 -53 24 -52
rect 24 -53 25 -52
rect 25 -53 26 -52
rect 40 -53 41 -52
rect 41 -53 42 -52
rect 42 -53 43 -52
rect 43 -53 44 -52
rect 44 -53 45 -52
rect 45 -53 46 -52
rect 46 -53 47 -52
rect 47 -53 48 -52
rect 48 -53 49 -52
rect 49 -53 50 -52
rect 50 -53 51 -52
rect 51 -53 52 -52
rect 52 -53 53 -52
rect 53 -53 54 -52
rect 54 -53 55 -52
rect 55 -53 56 -52
rect 56 -53 57 -52
rect 57 -53 58 -52
rect 72 -53 73 -52
rect 73 -53 74 -52
rect 74 -53 75 -52
rect 75 -53 76 -52
rect 76 -53 77 -52
rect 77 -53 78 -52
rect 78 -53 79 -52
rect 79 -53 80 -52
rect 80 -53 81 -52
rect 81 -53 82 -52
rect 82 -53 83 -52
rect 83 -53 84 -52
rect 84 -53 85 -52
rect 85 -53 86 -52
rect 86 -53 87 -52
rect 87 -53 88 -52
rect 88 -53 89 -52
rect 89 -53 90 -52
rect 104 -53 105 -52
rect 105 -53 106 -52
rect 106 -53 107 -52
rect 107 -53 108 -52
rect 108 -53 109 -52
rect 109 -53 110 -52
rect 110 -53 111 -52
rect 111 -53 112 -52
rect 112 -53 113 -52
rect 113 -53 114 -52
rect 114 -53 115 -52
rect 115 -53 116 -52
rect 116 -53 117 -52
rect 117 -53 118 -52
rect 118 -53 119 -52
rect 119 -53 120 -52
rect 120 -53 121 -52
rect 121 -53 122 -52
rect 136 -53 137 -52
rect 137 -53 138 -52
rect 138 -53 139 -52
rect 139 -53 140 -52
rect 140 -53 141 -52
rect 141 -53 142 -52
rect 142 -53 143 -52
rect 143 -53 144 -52
rect 144 -53 145 -52
rect 145 -53 146 -52
rect 146 -53 147 -52
rect 147 -53 148 -52
rect 148 -53 149 -52
rect 149 -53 150 -52
rect 150 -53 151 -52
rect 151 -53 152 -52
rect 152 -53 153 -52
rect 153 -53 154 -52
rect 168 -53 169 -52
rect 169 -53 170 -52
rect 170 -53 171 -52
rect 171 -53 172 -52
rect 172 -53 173 -52
rect 173 -53 174 -52
rect 174 -53 175 -52
rect 175 -53 176 -52
rect 176 -53 177 -52
rect 177 -53 178 -52
rect 178 -53 179 -52
rect 179 -53 180 -52
rect 180 -53 181 -52
rect 181 -53 182 -52
rect 182 -53 183 -52
rect 183 -53 184 -52
rect 184 -53 185 -52
rect 185 -53 186 -52
rect 186 -53 187 -52
rect 187 -53 188 -52
rect 188 -53 189 -52
rect 189 -53 190 -52
rect 190 -53 191 -52
rect 191 -53 192 -52
rect 192 -53 193 -52
rect 193 -53 194 -52
rect 194 -53 195 -52
rect 195 -53 196 -52
rect 196 -53 197 -52
rect 197 -53 198 -52
rect 198 -53 199 -52
rect 199 -53 200 -52
rect 200 -53 201 -52
rect 201 -53 202 -52
rect 202 -53 203 -52
rect 203 -53 204 -52
rect 204 -53 205 -52
rect 205 -53 206 -52
rect 206 -53 207 -52
rect 207 -53 208 -52
rect 208 -53 209 -52
rect 209 -53 210 -52
rect 210 -53 211 -52
rect 211 -53 212 -52
rect 212 -53 213 -52
rect 213 -53 214 -52
rect 214 -53 215 -52
rect 215 -53 216 -52
rect 216 -53 217 -52
rect 217 -53 218 -52
rect 218 -53 219 -52
rect 219 -53 220 -52
rect 220 -53 221 -52
rect 221 -53 222 -52
rect 222 -53 223 -52
rect 223 -53 224 -52
rect 224 -53 225 -52
rect 225 -53 226 -52
rect 226 -53 227 -52
rect 227 -53 228 -52
rect 228 -53 229 -52
rect 229 -53 230 -52
rect 230 -53 231 -52
rect 231 -53 232 -52
rect 232 -53 233 -52
rect 233 -53 234 -52
rect 234 -53 235 -52
rect 235 -53 236 -52
rect 236 -53 237 -52
rect 237 -53 238 -52
rect 238 -53 239 -52
rect 239 -53 240 -52
rect 240 -53 241 -52
rect 241 -53 242 -52
rect 242 -53 243 -52
rect 243 -53 244 -52
rect 244 -53 245 -52
rect 245 -53 246 -52
rect 246 -53 247 -52
rect 247 -53 248 -52
rect 248 -53 249 -52
rect 249 -53 250 -52
rect 250 -53 251 -52
rect 251 -53 252 -52
rect 252 -53 253 -52
rect 253 -53 254 -52
rect 254 -53 255 -52
rect 255 -53 256 -52
rect 256 -53 257 -52
rect 257 -53 258 -52
rect 258 -53 259 -52
rect 259 -53 260 -52
rect 260 -53 261 -52
rect 261 -53 262 -52
rect 262 -53 263 -52
rect 263 -53 264 -52
rect 264 -53 265 -52
rect 265 -53 266 -52
rect 266 -53 267 -52
rect 267 -53 268 -52
rect 268 -53 269 -52
rect 269 -53 270 -52
rect 270 -53 271 -52
rect 271 -53 272 -52
rect 272 -53 273 -52
rect 273 -53 274 -52
rect 274 -53 275 -52
rect 275 -53 276 -52
rect 276 -53 277 -52
rect 277 -53 278 -52
rect 278 -53 279 -52
rect 279 -53 280 -52
rect 280 -53 281 -52
rect 281 -53 282 -52
rect 282 -53 283 -52
rect 283 -53 284 -52
rect 284 -53 285 -52
rect 285 -53 286 -52
rect 286 -53 287 -52
rect 287 -53 288 -52
rect 288 -53 289 -52
rect 289 -53 290 -52
rect 290 -53 291 -52
rect 291 -53 292 -52
rect 292 -53 293 -52
rect 293 -53 294 -52
rect 294 -53 295 -52
rect 295 -53 296 -52
rect 296 -53 297 -52
rect 297 -53 298 -52
rect 298 -53 299 -52
rect 299 -53 300 -52
rect 300 -53 301 -52
rect 301 -53 302 -52
rect 302 -53 303 -52
rect 303 -53 304 -52
rect 304 -53 305 -52
rect 305 -53 306 -52
rect 306 -53 307 -52
rect 307 -53 308 -52
rect 308 -53 309 -52
rect 309 -53 310 -52
rect 310 -53 311 -52
rect 311 -53 312 -52
rect 312 -53 313 -52
rect 313 -53 314 -52
rect 314 -53 315 -52
rect 315 -53 316 -52
rect 316 -53 317 -52
rect 317 -53 318 -52
rect 318 -53 319 -52
rect 319 -53 320 -52
rect 320 -53 321 -52
rect 321 -53 322 -52
rect 322 -53 323 -52
rect 323 -53 324 -52
rect 324 -53 325 -52
rect 325 -53 326 -52
rect 326 -53 327 -52
rect 327 -53 328 -52
rect 328 -53 329 -52
rect 329 -53 330 -52
rect 330 -53 331 -52
rect 331 -53 332 -52
rect 332 -53 333 -52
rect 333 -53 334 -52
rect 334 -53 335 -52
rect 335 -53 336 -52
rect 336 -53 337 -52
rect 337 -53 338 -52
rect 338 -53 339 -52
rect 339 -53 340 -52
rect 340 -53 341 -52
rect 341 -53 342 -52
rect 342 -53 343 -52
rect 343 -53 344 -52
rect 344 -53 345 -52
rect 345 -53 346 -52
rect 346 -53 347 -52
rect 347 -53 348 -52
rect 348 -53 349 -52
rect 349 -53 350 -52
rect 350 -53 351 -52
rect 351 -53 352 -52
rect 352 -53 353 -52
rect 353 -53 354 -52
rect 354 -53 355 -52
rect 355 -53 356 -52
rect 356 -53 357 -52
rect 357 -53 358 -52
rect 358 -53 359 -52
rect 359 -53 360 -52
rect 360 -53 361 -52
rect 361 -53 362 -52
rect 362 -53 363 -52
rect 363 -53 364 -52
rect 364 -53 365 -52
rect 365 -53 366 -52
rect 366 -53 367 -52
rect 367 -53 368 -52
rect 368 -53 369 -52
rect 369 -53 370 -52
rect 370 -53 371 -52
rect 371 -53 372 -52
rect 372 -53 373 -52
rect 373 -53 374 -52
rect 374 -53 375 -52
rect 375 -53 376 -52
rect 376 -53 377 -52
rect 377 -53 378 -52
rect 378 -53 379 -52
rect 379 -53 380 -52
rect 380 -53 381 -52
rect 381 -53 382 -52
rect 382 -53 383 -52
rect 383 -53 384 -52
rect 384 -53 385 -52
rect 385 -53 386 -52
rect 386 -53 387 -52
rect 387 -53 388 -52
rect 388 -53 389 -52
rect 389 -53 390 -52
rect 390 -53 391 -52
rect 391 -53 392 -52
rect 392 -53 393 -52
rect 393 -53 394 -52
rect 394 -53 395 -52
rect 395 -53 396 -52
rect 396 -53 397 -52
rect 397 -53 398 -52
rect 398 -53 399 -52
rect 399 -53 400 -52
rect 400 -53 401 -52
rect 401 -53 402 -52
rect 402 -53 403 -52
rect 403 -53 404 -52
rect 404 -53 405 -52
rect 405 -53 406 -52
rect 406 -53 407 -52
rect 407 -53 408 -52
rect 408 -53 409 -52
rect 409 -53 410 -52
rect 410 -53 411 -52
rect 411 -53 412 -52
rect 412 -53 413 -52
rect 413 -53 414 -52
rect 414 -53 415 -52
rect 415 -53 416 -52
rect 416 -53 417 -52
rect 417 -53 418 -52
rect 418 -53 419 -52
rect 419 -53 420 -52
rect 420 -53 421 -52
rect 421 -53 422 -52
rect 422 -53 423 -52
rect 423 -53 424 -52
rect 424 -53 425 -52
rect 425 -53 426 -52
rect 426 -53 427 -52
rect 427 -53 428 -52
rect 428 -53 429 -52
rect 429 -53 430 -52
rect 430 -53 431 -52
rect 431 -53 432 -52
rect 432 -53 433 -52
rect 433 -53 434 -52
rect 434 -53 435 -52
rect 435 -53 436 -52
rect 436 -53 437 -52
rect 437 -53 438 -52
rect 438 -53 439 -52
rect 439 -53 440 -52
rect 440 -53 441 -52
rect 441 -53 442 -52
rect 442 -53 443 -52
rect 443 -53 444 -52
rect 444 -53 445 -52
rect 445 -53 446 -52
rect 446 -53 447 -52
rect 447 -53 448 -52
rect 448 -53 449 -52
rect 449 -53 450 -52
rect 450 -53 451 -52
rect 451 -53 452 -52
rect 452 -53 453 -52
rect 453 -53 454 -52
rect 454 -53 455 -52
rect 455 -53 456 -52
rect 456 -53 457 -52
rect 457 -53 458 -52
rect 458 -53 459 -52
rect 459 -53 460 -52
rect 460 -53 461 -52
rect 461 -53 462 -52
rect 462 -53 463 -52
rect 463 -53 464 -52
rect 464 -53 465 -52
rect 465 -53 466 -52
rect 466 -53 467 -52
rect 467 -53 468 -52
rect 468 -53 469 -52
rect 469 -53 470 -52
rect 470 -53 471 -52
rect 471 -53 472 -52
rect 472 -53 473 -52
rect 473 -53 474 -52
rect 474 -53 475 -52
rect 475 -53 476 -52
rect 476 -53 477 -52
rect 477 -53 478 -52
rect 478 -53 479 -52
rect 479 -53 480 -52
rect 2 -54 3 -53
rect 3 -54 4 -53
rect 4 -54 5 -53
rect 5 -54 6 -53
rect 6 -54 7 -53
rect 7 -54 8 -53
rect 8 -54 9 -53
rect 9 -54 10 -53
rect 10 -54 11 -53
rect 11 -54 12 -53
rect 12 -54 13 -53
rect 13 -54 14 -53
rect 14 -54 15 -53
rect 15 -54 16 -53
rect 16 -54 17 -53
rect 17 -54 18 -53
rect 18 -54 19 -53
rect 19 -54 20 -53
rect 20 -54 21 -53
rect 21 -54 22 -53
rect 22 -54 23 -53
rect 23 -54 24 -53
rect 24 -54 25 -53
rect 25 -54 26 -53
rect 26 -54 27 -53
rect 39 -54 40 -53
rect 40 -54 41 -53
rect 41 -54 42 -53
rect 42 -54 43 -53
rect 43 -54 44 -53
rect 44 -54 45 -53
rect 45 -54 46 -53
rect 46 -54 47 -53
rect 47 -54 48 -53
rect 48 -54 49 -53
rect 49 -54 50 -53
rect 50 -54 51 -53
rect 51 -54 52 -53
rect 52 -54 53 -53
rect 53 -54 54 -53
rect 54 -54 55 -53
rect 55 -54 56 -53
rect 56 -54 57 -53
rect 57 -54 58 -53
rect 58 -54 59 -53
rect 71 -54 72 -53
rect 72 -54 73 -53
rect 73 -54 74 -53
rect 74 -54 75 -53
rect 75 -54 76 -53
rect 76 -54 77 -53
rect 77 -54 78 -53
rect 78 -54 79 -53
rect 79 -54 80 -53
rect 80 -54 81 -53
rect 81 -54 82 -53
rect 82 -54 83 -53
rect 83 -54 84 -53
rect 84 -54 85 -53
rect 85 -54 86 -53
rect 86 -54 87 -53
rect 87 -54 88 -53
rect 88 -54 89 -53
rect 89 -54 90 -53
rect 90 -54 91 -53
rect 103 -54 104 -53
rect 104 -54 105 -53
rect 105 -54 106 -53
rect 106 -54 107 -53
rect 107 -54 108 -53
rect 108 -54 109 -53
rect 109 -54 110 -53
rect 110 -54 111 -53
rect 111 -54 112 -53
rect 112 -54 113 -53
rect 113 -54 114 -53
rect 114 -54 115 -53
rect 115 -54 116 -53
rect 116 -54 117 -53
rect 117 -54 118 -53
rect 118 -54 119 -53
rect 119 -54 120 -53
rect 120 -54 121 -53
rect 121 -54 122 -53
rect 122 -54 123 -53
rect 135 -54 136 -53
rect 136 -54 137 -53
rect 137 -54 138 -53
rect 138 -54 139 -53
rect 139 -54 140 -53
rect 140 -54 141 -53
rect 141 -54 142 -53
rect 142 -54 143 -53
rect 143 -54 144 -53
rect 144 -54 145 -53
rect 145 -54 146 -53
rect 146 -54 147 -53
rect 147 -54 148 -53
rect 148 -54 149 -53
rect 149 -54 150 -53
rect 150 -54 151 -53
rect 151 -54 152 -53
rect 152 -54 153 -53
rect 153 -54 154 -53
rect 154 -54 155 -53
rect 167 -54 168 -53
rect 168 -54 169 -53
rect 169 -54 170 -53
rect 170 -54 171 -53
rect 171 -54 172 -53
rect 172 -54 173 -53
rect 173 -54 174 -53
rect 174 -54 175 -53
rect 175 -54 176 -53
rect 176 -54 177 -53
rect 177 -54 178 -53
rect 178 -54 179 -53
rect 179 -54 180 -53
rect 180 -54 181 -53
rect 181 -54 182 -53
rect 182 -54 183 -53
rect 183 -54 184 -53
rect 184 -54 185 -53
rect 185 -54 186 -53
rect 186 -54 187 -53
rect 187 -54 188 -53
rect 188 -54 189 -53
rect 189 -54 190 -53
rect 190 -54 191 -53
rect 191 -54 192 -53
rect 192 -54 193 -53
rect 193 -54 194 -53
rect 194 -54 195 -53
rect 195 -54 196 -53
rect 196 -54 197 -53
rect 197 -54 198 -53
rect 198 -54 199 -53
rect 199 -54 200 -53
rect 200 -54 201 -53
rect 201 -54 202 -53
rect 202 -54 203 -53
rect 203 -54 204 -53
rect 204 -54 205 -53
rect 205 -54 206 -53
rect 206 -54 207 -53
rect 207 -54 208 -53
rect 208 -54 209 -53
rect 209 -54 210 -53
rect 210 -54 211 -53
rect 211 -54 212 -53
rect 212 -54 213 -53
rect 213 -54 214 -53
rect 214 -54 215 -53
rect 215 -54 216 -53
rect 216 -54 217 -53
rect 217 -54 218 -53
rect 218 -54 219 -53
rect 219 -54 220 -53
rect 220 -54 221 -53
rect 221 -54 222 -53
rect 222 -54 223 -53
rect 223 -54 224 -53
rect 224 -54 225 -53
rect 225 -54 226 -53
rect 226 -54 227 -53
rect 227 -54 228 -53
rect 228 -54 229 -53
rect 229 -54 230 -53
rect 230 -54 231 -53
rect 231 -54 232 -53
rect 232 -54 233 -53
rect 233 -54 234 -53
rect 234 -54 235 -53
rect 235 -54 236 -53
rect 236 -54 237 -53
rect 237 -54 238 -53
rect 238 -54 239 -53
rect 239 -54 240 -53
rect 240 -54 241 -53
rect 241 -54 242 -53
rect 242 -54 243 -53
rect 243 -54 244 -53
rect 244 -54 245 -53
rect 245 -54 246 -53
rect 246 -54 247 -53
rect 247 -54 248 -53
rect 248 -54 249 -53
rect 249 -54 250 -53
rect 250 -54 251 -53
rect 251 -54 252 -53
rect 252 -54 253 -53
rect 253 -54 254 -53
rect 254 -54 255 -53
rect 255 -54 256 -53
rect 256 -54 257 -53
rect 257 -54 258 -53
rect 258 -54 259 -53
rect 259 -54 260 -53
rect 260 -54 261 -53
rect 261 -54 262 -53
rect 262 -54 263 -53
rect 263 -54 264 -53
rect 264 -54 265 -53
rect 265 -54 266 -53
rect 266 -54 267 -53
rect 267 -54 268 -53
rect 268 -54 269 -53
rect 269 -54 270 -53
rect 270 -54 271 -53
rect 271 -54 272 -53
rect 272 -54 273 -53
rect 273 -54 274 -53
rect 274 -54 275 -53
rect 275 -54 276 -53
rect 276 -54 277 -53
rect 277 -54 278 -53
rect 278 -54 279 -53
rect 279 -54 280 -53
rect 280 -54 281 -53
rect 281 -54 282 -53
rect 282 -54 283 -53
rect 283 -54 284 -53
rect 284 -54 285 -53
rect 285 -54 286 -53
rect 286 -54 287 -53
rect 287 -54 288 -53
rect 288 -54 289 -53
rect 289 -54 290 -53
rect 290 -54 291 -53
rect 291 -54 292 -53
rect 292 -54 293 -53
rect 293 -54 294 -53
rect 294 -54 295 -53
rect 295 -54 296 -53
rect 296 -54 297 -53
rect 297 -54 298 -53
rect 298 -54 299 -53
rect 299 -54 300 -53
rect 300 -54 301 -53
rect 301 -54 302 -53
rect 302 -54 303 -53
rect 303 -54 304 -53
rect 304 -54 305 -53
rect 305 -54 306 -53
rect 306 -54 307 -53
rect 307 -54 308 -53
rect 308 -54 309 -53
rect 309 -54 310 -53
rect 310 -54 311 -53
rect 311 -54 312 -53
rect 312 -54 313 -53
rect 313 -54 314 -53
rect 314 -54 315 -53
rect 315 -54 316 -53
rect 316 -54 317 -53
rect 317 -54 318 -53
rect 318 -54 319 -53
rect 319 -54 320 -53
rect 320 -54 321 -53
rect 321 -54 322 -53
rect 322 -54 323 -53
rect 323 -54 324 -53
rect 324 -54 325 -53
rect 325 -54 326 -53
rect 326 -54 327 -53
rect 327 -54 328 -53
rect 328 -54 329 -53
rect 329 -54 330 -53
rect 330 -54 331 -53
rect 331 -54 332 -53
rect 332 -54 333 -53
rect 333 -54 334 -53
rect 334 -54 335 -53
rect 335 -54 336 -53
rect 336 -54 337 -53
rect 337 -54 338 -53
rect 338 -54 339 -53
rect 339 -54 340 -53
rect 340 -54 341 -53
rect 341 -54 342 -53
rect 342 -54 343 -53
rect 343 -54 344 -53
rect 344 -54 345 -53
rect 345 -54 346 -53
rect 346 -54 347 -53
rect 347 -54 348 -53
rect 348 -54 349 -53
rect 349 -54 350 -53
rect 350 -54 351 -53
rect 351 -54 352 -53
rect 352 -54 353 -53
rect 353 -54 354 -53
rect 354 -54 355 -53
rect 355 -54 356 -53
rect 356 -54 357 -53
rect 357 -54 358 -53
rect 358 -54 359 -53
rect 359 -54 360 -53
rect 360 -54 361 -53
rect 361 -54 362 -53
rect 362 -54 363 -53
rect 363 -54 364 -53
rect 364 -54 365 -53
rect 365 -54 366 -53
rect 366 -54 367 -53
rect 367 -54 368 -53
rect 368 -54 369 -53
rect 369 -54 370 -53
rect 370 -54 371 -53
rect 371 -54 372 -53
rect 372 -54 373 -53
rect 373 -54 374 -53
rect 374 -54 375 -53
rect 375 -54 376 -53
rect 376 -54 377 -53
rect 377 -54 378 -53
rect 378 -54 379 -53
rect 379 -54 380 -53
rect 380 -54 381 -53
rect 381 -54 382 -53
rect 382 -54 383 -53
rect 383 -54 384 -53
rect 384 -54 385 -53
rect 385 -54 386 -53
rect 386 -54 387 -53
rect 387 -54 388 -53
rect 388 -54 389 -53
rect 389 -54 390 -53
rect 390 -54 391 -53
rect 391 -54 392 -53
rect 392 -54 393 -53
rect 393 -54 394 -53
rect 394 -54 395 -53
rect 395 -54 396 -53
rect 396 -54 397 -53
rect 397 -54 398 -53
rect 398 -54 399 -53
rect 399 -54 400 -53
rect 400 -54 401 -53
rect 401 -54 402 -53
rect 402 -54 403 -53
rect 403 -54 404 -53
rect 404 -54 405 -53
rect 405 -54 406 -53
rect 406 -54 407 -53
rect 407 -54 408 -53
rect 408 -54 409 -53
rect 409 -54 410 -53
rect 410 -54 411 -53
rect 411 -54 412 -53
rect 412 -54 413 -53
rect 413 -54 414 -53
rect 414 -54 415 -53
rect 415 -54 416 -53
rect 416 -54 417 -53
rect 417 -54 418 -53
rect 418 -54 419 -53
rect 419 -54 420 -53
rect 420 -54 421 -53
rect 421 -54 422 -53
rect 422 -54 423 -53
rect 423 -54 424 -53
rect 424 -54 425 -53
rect 425 -54 426 -53
rect 426 -54 427 -53
rect 427 -54 428 -53
rect 428 -54 429 -53
rect 429 -54 430 -53
rect 430 -54 431 -53
rect 431 -54 432 -53
rect 432 -54 433 -53
rect 433 -54 434 -53
rect 434 -54 435 -53
rect 435 -54 436 -53
rect 436 -54 437 -53
rect 437 -54 438 -53
rect 438 -54 439 -53
rect 439 -54 440 -53
rect 440 -54 441 -53
rect 441 -54 442 -53
rect 442 -54 443 -53
rect 443 -54 444 -53
rect 444 -54 445 -53
rect 445 -54 446 -53
rect 446 -54 447 -53
rect 447 -54 448 -53
rect 448 -54 449 -53
rect 449 -54 450 -53
rect 450 -54 451 -53
rect 451 -54 452 -53
rect 452 -54 453 -53
rect 453 -54 454 -53
rect 454 -54 455 -53
rect 455 -54 456 -53
rect 456 -54 457 -53
rect 457 -54 458 -53
rect 458 -54 459 -53
rect 459 -54 460 -53
rect 460 -54 461 -53
rect 461 -54 462 -53
rect 462 -54 463 -53
rect 463 -54 464 -53
rect 464 -54 465 -53
rect 465 -54 466 -53
rect 466 -54 467 -53
rect 467 -54 468 -53
rect 468 -54 469 -53
rect 469 -54 470 -53
rect 470 -54 471 -53
rect 471 -54 472 -53
rect 472 -54 473 -53
rect 473 -54 474 -53
rect 474 -54 475 -53
rect 475 -54 476 -53
rect 476 -54 477 -53
rect 477 -54 478 -53
rect 478 -54 479 -53
rect 479 -54 480 -53
rect 2 -55 3 -54
rect 3 -55 4 -54
rect 4 -55 5 -54
rect 5 -55 6 -54
rect 6 -55 7 -54
rect 7 -55 8 -54
rect 8 -55 9 -54
rect 9 -55 10 -54
rect 10 -55 11 -54
rect 11 -55 12 -54
rect 12 -55 13 -54
rect 13 -55 14 -54
rect 14 -55 15 -54
rect 15 -55 16 -54
rect 16 -55 17 -54
rect 17 -55 18 -54
rect 18 -55 19 -54
rect 19 -55 20 -54
rect 20 -55 21 -54
rect 21 -55 22 -54
rect 22 -55 23 -54
rect 23 -55 24 -54
rect 24 -55 25 -54
rect 25 -55 26 -54
rect 26 -55 27 -54
rect 27 -55 28 -54
rect 38 -55 39 -54
rect 39 -55 40 -54
rect 40 -55 41 -54
rect 41 -55 42 -54
rect 42 -55 43 -54
rect 43 -55 44 -54
rect 44 -55 45 -54
rect 45 -55 46 -54
rect 46 -55 47 -54
rect 47 -55 48 -54
rect 48 -55 49 -54
rect 49 -55 50 -54
rect 50 -55 51 -54
rect 51 -55 52 -54
rect 52 -55 53 -54
rect 53 -55 54 -54
rect 54 -55 55 -54
rect 55 -55 56 -54
rect 56 -55 57 -54
rect 57 -55 58 -54
rect 58 -55 59 -54
rect 59 -55 60 -54
rect 70 -55 71 -54
rect 71 -55 72 -54
rect 72 -55 73 -54
rect 73 -55 74 -54
rect 74 -55 75 -54
rect 75 -55 76 -54
rect 76 -55 77 -54
rect 77 -55 78 -54
rect 78 -55 79 -54
rect 79 -55 80 -54
rect 80 -55 81 -54
rect 81 -55 82 -54
rect 82 -55 83 -54
rect 83 -55 84 -54
rect 84 -55 85 -54
rect 85 -55 86 -54
rect 86 -55 87 -54
rect 87 -55 88 -54
rect 88 -55 89 -54
rect 89 -55 90 -54
rect 90 -55 91 -54
rect 91 -55 92 -54
rect 102 -55 103 -54
rect 103 -55 104 -54
rect 104 -55 105 -54
rect 105 -55 106 -54
rect 106 -55 107 -54
rect 107 -55 108 -54
rect 108 -55 109 -54
rect 109 -55 110 -54
rect 110 -55 111 -54
rect 111 -55 112 -54
rect 112 -55 113 -54
rect 113 -55 114 -54
rect 114 -55 115 -54
rect 115 -55 116 -54
rect 116 -55 117 -54
rect 117 -55 118 -54
rect 118 -55 119 -54
rect 119 -55 120 -54
rect 120 -55 121 -54
rect 121 -55 122 -54
rect 122 -55 123 -54
rect 123 -55 124 -54
rect 134 -55 135 -54
rect 135 -55 136 -54
rect 136 -55 137 -54
rect 137 -55 138 -54
rect 138 -55 139 -54
rect 139 -55 140 -54
rect 140 -55 141 -54
rect 141 -55 142 -54
rect 142 -55 143 -54
rect 143 -55 144 -54
rect 144 -55 145 -54
rect 145 -55 146 -54
rect 146 -55 147 -54
rect 147 -55 148 -54
rect 148 -55 149 -54
rect 149 -55 150 -54
rect 150 -55 151 -54
rect 151 -55 152 -54
rect 152 -55 153 -54
rect 153 -55 154 -54
rect 154 -55 155 -54
rect 155 -55 156 -54
rect 166 -55 167 -54
rect 167 -55 168 -54
rect 168 -55 169 -54
rect 169 -55 170 -54
rect 170 -55 171 -54
rect 171 -55 172 -54
rect 172 -55 173 -54
rect 173 -55 174 -54
rect 174 -55 175 -54
rect 175 -55 176 -54
rect 176 -55 177 -54
rect 177 -55 178 -54
rect 178 -55 179 -54
rect 179 -55 180 -54
rect 180 -55 181 -54
rect 181 -55 182 -54
rect 182 -55 183 -54
rect 183 -55 184 -54
rect 184 -55 185 -54
rect 185 -55 186 -54
rect 186 -55 187 -54
rect 187 -55 188 -54
rect 188 -55 189 -54
rect 189 -55 190 -54
rect 190 -55 191 -54
rect 191 -55 192 -54
rect 192 -55 193 -54
rect 193 -55 194 -54
rect 194 -55 195 -54
rect 195 -55 196 -54
rect 196 -55 197 -54
rect 197 -55 198 -54
rect 198 -55 199 -54
rect 199 -55 200 -54
rect 200 -55 201 -54
rect 201 -55 202 -54
rect 202 -55 203 -54
rect 203 -55 204 -54
rect 204 -55 205 -54
rect 205 -55 206 -54
rect 206 -55 207 -54
rect 207 -55 208 -54
rect 208 -55 209 -54
rect 209 -55 210 -54
rect 210 -55 211 -54
rect 211 -55 212 -54
rect 212 -55 213 -54
rect 213 -55 214 -54
rect 214 -55 215 -54
rect 215 -55 216 -54
rect 216 -55 217 -54
rect 217 -55 218 -54
rect 218 -55 219 -54
rect 219 -55 220 -54
rect 220 -55 221 -54
rect 221 -55 222 -54
rect 222 -55 223 -54
rect 223 -55 224 -54
rect 224 -55 225 -54
rect 225 -55 226 -54
rect 226 -55 227 -54
rect 227 -55 228 -54
rect 228 -55 229 -54
rect 229 -55 230 -54
rect 230 -55 231 -54
rect 231 -55 232 -54
rect 232 -55 233 -54
rect 233 -55 234 -54
rect 234 -55 235 -54
rect 235 -55 236 -54
rect 236 -55 237 -54
rect 237 -55 238 -54
rect 238 -55 239 -54
rect 239 -55 240 -54
rect 240 -55 241 -54
rect 241 -55 242 -54
rect 242 -55 243 -54
rect 243 -55 244 -54
rect 244 -55 245 -54
rect 245 -55 246 -54
rect 246 -55 247 -54
rect 247 -55 248 -54
rect 248 -55 249 -54
rect 249 -55 250 -54
rect 250 -55 251 -54
rect 251 -55 252 -54
rect 252 -55 253 -54
rect 253 -55 254 -54
rect 254 -55 255 -54
rect 255 -55 256 -54
rect 256 -55 257 -54
rect 257 -55 258 -54
rect 258 -55 259 -54
rect 259 -55 260 -54
rect 260 -55 261 -54
rect 261 -55 262 -54
rect 262 -55 263 -54
rect 263 -55 264 -54
rect 264 -55 265 -54
rect 265 -55 266 -54
rect 266 -55 267 -54
rect 267 -55 268 -54
rect 268 -55 269 -54
rect 269 -55 270 -54
rect 270 -55 271 -54
rect 271 -55 272 -54
rect 272 -55 273 -54
rect 273 -55 274 -54
rect 274 -55 275 -54
rect 275 -55 276 -54
rect 276 -55 277 -54
rect 277 -55 278 -54
rect 278 -55 279 -54
rect 279 -55 280 -54
rect 280 -55 281 -54
rect 281 -55 282 -54
rect 282 -55 283 -54
rect 283 -55 284 -54
rect 284 -55 285 -54
rect 285 -55 286 -54
rect 286 -55 287 -54
rect 287 -55 288 -54
rect 288 -55 289 -54
rect 289 -55 290 -54
rect 290 -55 291 -54
rect 291 -55 292 -54
rect 292 -55 293 -54
rect 293 -55 294 -54
rect 294 -55 295 -54
rect 295 -55 296 -54
rect 296 -55 297 -54
rect 297 -55 298 -54
rect 298 -55 299 -54
rect 299 -55 300 -54
rect 300 -55 301 -54
rect 301 -55 302 -54
rect 302 -55 303 -54
rect 303 -55 304 -54
rect 304 -55 305 -54
rect 305 -55 306 -54
rect 306 -55 307 -54
rect 307 -55 308 -54
rect 308 -55 309 -54
rect 309 -55 310 -54
rect 310 -55 311 -54
rect 311 -55 312 -54
rect 312 -55 313 -54
rect 313 -55 314 -54
rect 314 -55 315 -54
rect 315 -55 316 -54
rect 316 -55 317 -54
rect 317 -55 318 -54
rect 318 -55 319 -54
rect 319 -55 320 -54
rect 320 -55 321 -54
rect 321 -55 322 -54
rect 322 -55 323 -54
rect 323 -55 324 -54
rect 324 -55 325 -54
rect 325 -55 326 -54
rect 326 -55 327 -54
rect 327 -55 328 -54
rect 328 -55 329 -54
rect 329 -55 330 -54
rect 330 -55 331 -54
rect 331 -55 332 -54
rect 332 -55 333 -54
rect 333 -55 334 -54
rect 334 -55 335 -54
rect 335 -55 336 -54
rect 336 -55 337 -54
rect 337 -55 338 -54
rect 338 -55 339 -54
rect 339 -55 340 -54
rect 340 -55 341 -54
rect 341 -55 342 -54
rect 342 -55 343 -54
rect 343 -55 344 -54
rect 344 -55 345 -54
rect 345 -55 346 -54
rect 346 -55 347 -54
rect 347 -55 348 -54
rect 348 -55 349 -54
rect 349 -55 350 -54
rect 350 -55 351 -54
rect 351 -55 352 -54
rect 352 -55 353 -54
rect 353 -55 354 -54
rect 354 -55 355 -54
rect 355 -55 356 -54
rect 356 -55 357 -54
rect 357 -55 358 -54
rect 358 -55 359 -54
rect 359 -55 360 -54
rect 360 -55 361 -54
rect 361 -55 362 -54
rect 362 -55 363 -54
rect 363 -55 364 -54
rect 364 -55 365 -54
rect 365 -55 366 -54
rect 366 -55 367 -54
rect 367 -55 368 -54
rect 368 -55 369 -54
rect 369 -55 370 -54
rect 370 -55 371 -54
rect 371 -55 372 -54
rect 372 -55 373 -54
rect 373 -55 374 -54
rect 374 -55 375 -54
rect 375 -55 376 -54
rect 376 -55 377 -54
rect 377 -55 378 -54
rect 378 -55 379 -54
rect 379 -55 380 -54
rect 380 -55 381 -54
rect 381 -55 382 -54
rect 382 -55 383 -54
rect 383 -55 384 -54
rect 384 -55 385 -54
rect 385 -55 386 -54
rect 386 -55 387 -54
rect 387 -55 388 -54
rect 388 -55 389 -54
rect 389 -55 390 -54
rect 390 -55 391 -54
rect 391 -55 392 -54
rect 392 -55 393 -54
rect 393 -55 394 -54
rect 394 -55 395 -54
rect 395 -55 396 -54
rect 396 -55 397 -54
rect 397 -55 398 -54
rect 398 -55 399 -54
rect 399 -55 400 -54
rect 400 -55 401 -54
rect 401 -55 402 -54
rect 402 -55 403 -54
rect 403 -55 404 -54
rect 404 -55 405 -54
rect 405 -55 406 -54
rect 406 -55 407 -54
rect 407 -55 408 -54
rect 408 -55 409 -54
rect 409 -55 410 -54
rect 410 -55 411 -54
rect 411 -55 412 -54
rect 412 -55 413 -54
rect 413 -55 414 -54
rect 414 -55 415 -54
rect 415 -55 416 -54
rect 416 -55 417 -54
rect 417 -55 418 -54
rect 418 -55 419 -54
rect 419 -55 420 -54
rect 420 -55 421 -54
rect 421 -55 422 -54
rect 422 -55 423 -54
rect 423 -55 424 -54
rect 424 -55 425 -54
rect 425 -55 426 -54
rect 426 -55 427 -54
rect 427 -55 428 -54
rect 428 -55 429 -54
rect 429 -55 430 -54
rect 430 -55 431 -54
rect 431 -55 432 -54
rect 432 -55 433 -54
rect 433 -55 434 -54
rect 434 -55 435 -54
rect 435 -55 436 -54
rect 436 -55 437 -54
rect 437 -55 438 -54
rect 438 -55 439 -54
rect 439 -55 440 -54
rect 440 -55 441 -54
rect 441 -55 442 -54
rect 442 -55 443 -54
rect 443 -55 444 -54
rect 444 -55 445 -54
rect 445 -55 446 -54
rect 446 -55 447 -54
rect 447 -55 448 -54
rect 448 -55 449 -54
rect 449 -55 450 -54
rect 450 -55 451 -54
rect 451 -55 452 -54
rect 452 -55 453 -54
rect 453 -55 454 -54
rect 454 -55 455 -54
rect 455 -55 456 -54
rect 456 -55 457 -54
rect 457 -55 458 -54
rect 458 -55 459 -54
rect 459 -55 460 -54
rect 460 -55 461 -54
rect 461 -55 462 -54
rect 462 -55 463 -54
rect 463 -55 464 -54
rect 464 -55 465 -54
rect 465 -55 466 -54
rect 466 -55 467 -54
rect 467 -55 468 -54
rect 468 -55 469 -54
rect 469 -55 470 -54
rect 470 -55 471 -54
rect 471 -55 472 -54
rect 472 -55 473 -54
rect 473 -55 474 -54
rect 474 -55 475 -54
rect 475 -55 476 -54
rect 476 -55 477 -54
rect 477 -55 478 -54
rect 478 -55 479 -54
rect 479 -55 480 -54
rect 2 -56 3 -55
rect 3 -56 4 -55
rect 4 -56 5 -55
rect 5 -56 6 -55
rect 6 -56 7 -55
rect 7 -56 8 -55
rect 8 -56 9 -55
rect 9 -56 10 -55
rect 10 -56 11 -55
rect 11 -56 12 -55
rect 12 -56 13 -55
rect 13 -56 14 -55
rect 14 -56 15 -55
rect 15 -56 16 -55
rect 16 -56 17 -55
rect 17 -56 18 -55
rect 18 -56 19 -55
rect 19 -56 20 -55
rect 20 -56 21 -55
rect 21 -56 22 -55
rect 22 -56 23 -55
rect 23 -56 24 -55
rect 24 -56 25 -55
rect 25 -56 26 -55
rect 26 -56 27 -55
rect 27 -56 28 -55
rect 37 -56 38 -55
rect 38 -56 39 -55
rect 39 -56 40 -55
rect 40 -56 41 -55
rect 41 -56 42 -55
rect 42 -56 43 -55
rect 43 -56 44 -55
rect 44 -56 45 -55
rect 45 -56 46 -55
rect 46 -56 47 -55
rect 47 -56 48 -55
rect 48 -56 49 -55
rect 49 -56 50 -55
rect 50 -56 51 -55
rect 51 -56 52 -55
rect 52 -56 53 -55
rect 53 -56 54 -55
rect 54 -56 55 -55
rect 55 -56 56 -55
rect 56 -56 57 -55
rect 57 -56 58 -55
rect 58 -56 59 -55
rect 59 -56 60 -55
rect 69 -56 70 -55
rect 70 -56 71 -55
rect 71 -56 72 -55
rect 72 -56 73 -55
rect 73 -56 74 -55
rect 74 -56 75 -55
rect 75 -56 76 -55
rect 76 -56 77 -55
rect 77 -56 78 -55
rect 78 -56 79 -55
rect 79 -56 80 -55
rect 80 -56 81 -55
rect 81 -56 82 -55
rect 82 -56 83 -55
rect 83 -56 84 -55
rect 84 -56 85 -55
rect 85 -56 86 -55
rect 86 -56 87 -55
rect 87 -56 88 -55
rect 88 -56 89 -55
rect 89 -56 90 -55
rect 90 -56 91 -55
rect 91 -56 92 -55
rect 101 -56 102 -55
rect 102 -56 103 -55
rect 103 -56 104 -55
rect 104 -56 105 -55
rect 105 -56 106 -55
rect 106 -56 107 -55
rect 107 -56 108 -55
rect 108 -56 109 -55
rect 109 -56 110 -55
rect 110 -56 111 -55
rect 111 -56 112 -55
rect 112 -56 113 -55
rect 113 -56 114 -55
rect 114 -56 115 -55
rect 115 -56 116 -55
rect 116 -56 117 -55
rect 117 -56 118 -55
rect 118 -56 119 -55
rect 119 -56 120 -55
rect 120 -56 121 -55
rect 121 -56 122 -55
rect 122 -56 123 -55
rect 123 -56 124 -55
rect 133 -56 134 -55
rect 134 -56 135 -55
rect 135 -56 136 -55
rect 136 -56 137 -55
rect 137 -56 138 -55
rect 138 -56 139 -55
rect 139 -56 140 -55
rect 140 -56 141 -55
rect 141 -56 142 -55
rect 142 -56 143 -55
rect 143 -56 144 -55
rect 144 -56 145 -55
rect 145 -56 146 -55
rect 146 -56 147 -55
rect 147 -56 148 -55
rect 148 -56 149 -55
rect 149 -56 150 -55
rect 150 -56 151 -55
rect 151 -56 152 -55
rect 152 -56 153 -55
rect 153 -56 154 -55
rect 154 -56 155 -55
rect 155 -56 156 -55
rect 165 -56 166 -55
rect 166 -56 167 -55
rect 167 -56 168 -55
rect 168 -56 169 -55
rect 169 -56 170 -55
rect 170 -56 171 -55
rect 171 -56 172 -55
rect 172 -56 173 -55
rect 173 -56 174 -55
rect 174 -56 175 -55
rect 175 -56 176 -55
rect 176 -56 177 -55
rect 177 -56 178 -55
rect 178 -56 179 -55
rect 179 -56 180 -55
rect 180 -56 181 -55
rect 181 -56 182 -55
rect 182 -56 183 -55
rect 183 -56 184 -55
rect 184 -56 185 -55
rect 185 -56 186 -55
rect 186 -56 187 -55
rect 187 -56 188 -55
rect 188 -56 189 -55
rect 189 -56 190 -55
rect 190 -56 191 -55
rect 191 -56 192 -55
rect 192 -56 193 -55
rect 193 -56 194 -55
rect 194 -56 195 -55
rect 195 -56 196 -55
rect 196 -56 197 -55
rect 197 -56 198 -55
rect 198 -56 199 -55
rect 199 -56 200 -55
rect 200 -56 201 -55
rect 201 -56 202 -55
rect 202 -56 203 -55
rect 203 -56 204 -55
rect 204 -56 205 -55
rect 205 -56 206 -55
rect 206 -56 207 -55
rect 207 -56 208 -55
rect 208 -56 209 -55
rect 209 -56 210 -55
rect 210 -56 211 -55
rect 211 -56 212 -55
rect 212 -56 213 -55
rect 213 -56 214 -55
rect 214 -56 215 -55
rect 215 -56 216 -55
rect 216 -56 217 -55
rect 217 -56 218 -55
rect 218 -56 219 -55
rect 219 -56 220 -55
rect 220 -56 221 -55
rect 221 -56 222 -55
rect 222 -56 223 -55
rect 223 -56 224 -55
rect 224 -56 225 -55
rect 225 -56 226 -55
rect 226 -56 227 -55
rect 227 -56 228 -55
rect 228 -56 229 -55
rect 229 -56 230 -55
rect 230 -56 231 -55
rect 231 -56 232 -55
rect 232 -56 233 -55
rect 233 -56 234 -55
rect 234 -56 235 -55
rect 235 -56 236 -55
rect 236 -56 237 -55
rect 237 -56 238 -55
rect 238 -56 239 -55
rect 239 -56 240 -55
rect 240 -56 241 -55
rect 241 -56 242 -55
rect 242 -56 243 -55
rect 243 -56 244 -55
rect 244 -56 245 -55
rect 245 -56 246 -55
rect 246 -56 247 -55
rect 247 -56 248 -55
rect 248 -56 249 -55
rect 249 -56 250 -55
rect 250 -56 251 -55
rect 251 -56 252 -55
rect 252 -56 253 -55
rect 253 -56 254 -55
rect 254 -56 255 -55
rect 255 -56 256 -55
rect 256 -56 257 -55
rect 257 -56 258 -55
rect 258 -56 259 -55
rect 259 -56 260 -55
rect 260 -56 261 -55
rect 261 -56 262 -55
rect 262 -56 263 -55
rect 263 -56 264 -55
rect 264 -56 265 -55
rect 265 -56 266 -55
rect 266 -56 267 -55
rect 267 -56 268 -55
rect 268 -56 269 -55
rect 269 -56 270 -55
rect 270 -56 271 -55
rect 271 -56 272 -55
rect 272 -56 273 -55
rect 273 -56 274 -55
rect 274 -56 275 -55
rect 275 -56 276 -55
rect 276 -56 277 -55
rect 277 -56 278 -55
rect 278 -56 279 -55
rect 279 -56 280 -55
rect 280 -56 281 -55
rect 281 -56 282 -55
rect 282 -56 283 -55
rect 283 -56 284 -55
rect 284 -56 285 -55
rect 285 -56 286 -55
rect 286 -56 287 -55
rect 287 -56 288 -55
rect 288 -56 289 -55
rect 289 -56 290 -55
rect 290 -56 291 -55
rect 291 -56 292 -55
rect 292 -56 293 -55
rect 293 -56 294 -55
rect 294 -56 295 -55
rect 295 -56 296 -55
rect 296 -56 297 -55
rect 297 -56 298 -55
rect 298 -56 299 -55
rect 299 -56 300 -55
rect 300 -56 301 -55
rect 301 -56 302 -55
rect 302 -56 303 -55
rect 303 -56 304 -55
rect 304 -56 305 -55
rect 305 -56 306 -55
rect 306 -56 307 -55
rect 307 -56 308 -55
rect 308 -56 309 -55
rect 309 -56 310 -55
rect 310 -56 311 -55
rect 311 -56 312 -55
rect 312 -56 313 -55
rect 313 -56 314 -55
rect 314 -56 315 -55
rect 315 -56 316 -55
rect 316 -56 317 -55
rect 317 -56 318 -55
rect 318 -56 319 -55
rect 319 -56 320 -55
rect 320 -56 321 -55
rect 321 -56 322 -55
rect 322 -56 323 -55
rect 323 -56 324 -55
rect 324 -56 325 -55
rect 325 -56 326 -55
rect 326 -56 327 -55
rect 327 -56 328 -55
rect 328 -56 329 -55
rect 329 -56 330 -55
rect 330 -56 331 -55
rect 331 -56 332 -55
rect 332 -56 333 -55
rect 333 -56 334 -55
rect 334 -56 335 -55
rect 335 -56 336 -55
rect 336 -56 337 -55
rect 337 -56 338 -55
rect 338 -56 339 -55
rect 339 -56 340 -55
rect 340 -56 341 -55
rect 341 -56 342 -55
rect 342 -56 343 -55
rect 343 -56 344 -55
rect 344 -56 345 -55
rect 345 -56 346 -55
rect 346 -56 347 -55
rect 347 -56 348 -55
rect 348 -56 349 -55
rect 349 -56 350 -55
rect 350 -56 351 -55
rect 351 -56 352 -55
rect 352 -56 353 -55
rect 353 -56 354 -55
rect 354 -56 355 -55
rect 355 -56 356 -55
rect 356 -56 357 -55
rect 357 -56 358 -55
rect 358 -56 359 -55
rect 359 -56 360 -55
rect 360 -56 361 -55
rect 361 -56 362 -55
rect 362 -56 363 -55
rect 363 -56 364 -55
rect 364 -56 365 -55
rect 365 -56 366 -55
rect 366 -56 367 -55
rect 367 -56 368 -55
rect 368 -56 369 -55
rect 369 -56 370 -55
rect 370 -56 371 -55
rect 371 -56 372 -55
rect 372 -56 373 -55
rect 373 -56 374 -55
rect 374 -56 375 -55
rect 375 -56 376 -55
rect 376 -56 377 -55
rect 377 -56 378 -55
rect 378 -56 379 -55
rect 379 -56 380 -55
rect 380 -56 381 -55
rect 381 -56 382 -55
rect 382 -56 383 -55
rect 383 -56 384 -55
rect 384 -56 385 -55
rect 385 -56 386 -55
rect 386 -56 387 -55
rect 387 -56 388 -55
rect 388 -56 389 -55
rect 389 -56 390 -55
rect 390 -56 391 -55
rect 391 -56 392 -55
rect 392 -56 393 -55
rect 393 -56 394 -55
rect 394 -56 395 -55
rect 395 -56 396 -55
rect 396 -56 397 -55
rect 397 -56 398 -55
rect 398 -56 399 -55
rect 399 -56 400 -55
rect 400 -56 401 -55
rect 401 -56 402 -55
rect 402 -56 403 -55
rect 403 -56 404 -55
rect 404 -56 405 -55
rect 405 -56 406 -55
rect 406 -56 407 -55
rect 407 -56 408 -55
rect 408 -56 409 -55
rect 409 -56 410 -55
rect 410 -56 411 -55
rect 411 -56 412 -55
rect 412 -56 413 -55
rect 413 -56 414 -55
rect 414 -56 415 -55
rect 415 -56 416 -55
rect 416 -56 417 -55
rect 417 -56 418 -55
rect 418 -56 419 -55
rect 419 -56 420 -55
rect 420 -56 421 -55
rect 421 -56 422 -55
rect 422 -56 423 -55
rect 423 -56 424 -55
rect 424 -56 425 -55
rect 425 -56 426 -55
rect 426 -56 427 -55
rect 427 -56 428 -55
rect 428 -56 429 -55
rect 429 -56 430 -55
rect 430 -56 431 -55
rect 431 -56 432 -55
rect 432 -56 433 -55
rect 433 -56 434 -55
rect 434 -56 435 -55
rect 435 -56 436 -55
rect 436 -56 437 -55
rect 437 -56 438 -55
rect 438 -56 439 -55
rect 439 -56 440 -55
rect 440 -56 441 -55
rect 441 -56 442 -55
rect 442 -56 443 -55
rect 443 -56 444 -55
rect 444 -56 445 -55
rect 445 -56 446 -55
rect 446 -56 447 -55
rect 447 -56 448 -55
rect 448 -56 449 -55
rect 449 -56 450 -55
rect 450 -56 451 -55
rect 451 -56 452 -55
rect 452 -56 453 -55
rect 453 -56 454 -55
rect 454 -56 455 -55
rect 455 -56 456 -55
rect 456 -56 457 -55
rect 457 -56 458 -55
rect 458 -56 459 -55
rect 459 -56 460 -55
rect 460 -56 461 -55
rect 461 -56 462 -55
rect 462 -56 463 -55
rect 463 -56 464 -55
rect 464 -56 465 -55
rect 465 -56 466 -55
rect 466 -56 467 -55
rect 467 -56 468 -55
rect 468 -56 469 -55
rect 469 -56 470 -55
rect 470 -56 471 -55
rect 471 -56 472 -55
rect 472 -56 473 -55
rect 473 -56 474 -55
rect 474 -56 475 -55
rect 475 -56 476 -55
rect 476 -56 477 -55
rect 477 -56 478 -55
rect 478 -56 479 -55
rect 479 -56 480 -55
rect 2 -57 3 -56
rect 3 -57 4 -56
rect 4 -57 5 -56
rect 5 -57 6 -56
rect 6 -57 7 -56
rect 7 -57 8 -56
rect 8 -57 9 -56
rect 9 -57 10 -56
rect 10 -57 11 -56
rect 11 -57 12 -56
rect 12 -57 13 -56
rect 13 -57 14 -56
rect 14 -57 15 -56
rect 15 -57 16 -56
rect 16 -57 17 -56
rect 17 -57 18 -56
rect 18 -57 19 -56
rect 19 -57 20 -56
rect 20 -57 21 -56
rect 21 -57 22 -56
rect 22 -57 23 -56
rect 23 -57 24 -56
rect 24 -57 25 -56
rect 25 -57 26 -56
rect 26 -57 27 -56
rect 27 -57 28 -56
rect 37 -57 38 -56
rect 38 -57 39 -56
rect 39 -57 40 -56
rect 40 -57 41 -56
rect 41 -57 42 -56
rect 42 -57 43 -56
rect 43 -57 44 -56
rect 44 -57 45 -56
rect 45 -57 46 -56
rect 46 -57 47 -56
rect 47 -57 48 -56
rect 48 -57 49 -56
rect 49 -57 50 -56
rect 50 -57 51 -56
rect 51 -57 52 -56
rect 52 -57 53 -56
rect 53 -57 54 -56
rect 54 -57 55 -56
rect 55 -57 56 -56
rect 56 -57 57 -56
rect 57 -57 58 -56
rect 58 -57 59 -56
rect 59 -57 60 -56
rect 69 -57 70 -56
rect 70 -57 71 -56
rect 71 -57 72 -56
rect 72 -57 73 -56
rect 73 -57 74 -56
rect 74 -57 75 -56
rect 75 -57 76 -56
rect 76 -57 77 -56
rect 77 -57 78 -56
rect 78 -57 79 -56
rect 79 -57 80 -56
rect 80 -57 81 -56
rect 81 -57 82 -56
rect 82 -57 83 -56
rect 83 -57 84 -56
rect 84 -57 85 -56
rect 85 -57 86 -56
rect 86 -57 87 -56
rect 87 -57 88 -56
rect 88 -57 89 -56
rect 89 -57 90 -56
rect 90 -57 91 -56
rect 91 -57 92 -56
rect 101 -57 102 -56
rect 102 -57 103 -56
rect 103 -57 104 -56
rect 104 -57 105 -56
rect 105 -57 106 -56
rect 106 -57 107 -56
rect 107 -57 108 -56
rect 108 -57 109 -56
rect 109 -57 110 -56
rect 110 -57 111 -56
rect 111 -57 112 -56
rect 112 -57 113 -56
rect 113 -57 114 -56
rect 114 -57 115 -56
rect 115 -57 116 -56
rect 116 -57 117 -56
rect 117 -57 118 -56
rect 118 -57 119 -56
rect 119 -57 120 -56
rect 120 -57 121 -56
rect 121 -57 122 -56
rect 122 -57 123 -56
rect 123 -57 124 -56
rect 133 -57 134 -56
rect 134 -57 135 -56
rect 135 -57 136 -56
rect 136 -57 137 -56
rect 137 -57 138 -56
rect 138 -57 139 -56
rect 139 -57 140 -56
rect 140 -57 141 -56
rect 141 -57 142 -56
rect 142 -57 143 -56
rect 143 -57 144 -56
rect 144 -57 145 -56
rect 145 -57 146 -56
rect 146 -57 147 -56
rect 147 -57 148 -56
rect 148 -57 149 -56
rect 149 -57 150 -56
rect 150 -57 151 -56
rect 151 -57 152 -56
rect 152 -57 153 -56
rect 153 -57 154 -56
rect 154 -57 155 -56
rect 155 -57 156 -56
rect 165 -57 166 -56
rect 166 -57 167 -56
rect 167 -57 168 -56
rect 168 -57 169 -56
rect 169 -57 170 -56
rect 170 -57 171 -56
rect 171 -57 172 -56
rect 172 -57 173 -56
rect 173 -57 174 -56
rect 174 -57 175 -56
rect 175 -57 176 -56
rect 176 -57 177 -56
rect 177 -57 178 -56
rect 178 -57 179 -56
rect 179 -57 180 -56
rect 180 -57 181 -56
rect 181 -57 182 -56
rect 182 -57 183 -56
rect 183 -57 184 -56
rect 184 -57 185 -56
rect 185 -57 186 -56
rect 186 -57 187 -56
rect 187 -57 188 -56
rect 188 -57 189 -56
rect 189 -57 190 -56
rect 190 -57 191 -56
rect 191 -57 192 -56
rect 192 -57 193 -56
rect 193 -57 194 -56
rect 194 -57 195 -56
rect 195 -57 196 -56
rect 196 -57 197 -56
rect 197 -57 198 -56
rect 198 -57 199 -56
rect 199 -57 200 -56
rect 200 -57 201 -56
rect 201 -57 202 -56
rect 202 -57 203 -56
rect 203 -57 204 -56
rect 204 -57 205 -56
rect 205 -57 206 -56
rect 206 -57 207 -56
rect 207 -57 208 -56
rect 208 -57 209 -56
rect 209 -57 210 -56
rect 210 -57 211 -56
rect 211 -57 212 -56
rect 212 -57 213 -56
rect 213 -57 214 -56
rect 214 -57 215 -56
rect 215 -57 216 -56
rect 216 -57 217 -56
rect 217 -57 218 -56
rect 218 -57 219 -56
rect 219 -57 220 -56
rect 220 -57 221 -56
rect 221 -57 222 -56
rect 222 -57 223 -56
rect 223 -57 224 -56
rect 224 -57 225 -56
rect 225 -57 226 -56
rect 226 -57 227 -56
rect 227 -57 228 -56
rect 228 -57 229 -56
rect 229 -57 230 -56
rect 230 -57 231 -56
rect 231 -57 232 -56
rect 232 -57 233 -56
rect 233 -57 234 -56
rect 234 -57 235 -56
rect 235 -57 236 -56
rect 236 -57 237 -56
rect 237 -57 238 -56
rect 238 -57 239 -56
rect 239 -57 240 -56
rect 240 -57 241 -56
rect 241 -57 242 -56
rect 242 -57 243 -56
rect 243 -57 244 -56
rect 244 -57 245 -56
rect 245 -57 246 -56
rect 246 -57 247 -56
rect 247 -57 248 -56
rect 248 -57 249 -56
rect 249 -57 250 -56
rect 250 -57 251 -56
rect 251 -57 252 -56
rect 252 -57 253 -56
rect 253 -57 254 -56
rect 254 -57 255 -56
rect 255 -57 256 -56
rect 256 -57 257 -56
rect 257 -57 258 -56
rect 258 -57 259 -56
rect 259 -57 260 -56
rect 260 -57 261 -56
rect 261 -57 262 -56
rect 262 -57 263 -56
rect 263 -57 264 -56
rect 264 -57 265 -56
rect 265 -57 266 -56
rect 266 -57 267 -56
rect 267 -57 268 -56
rect 268 -57 269 -56
rect 269 -57 270 -56
rect 270 -57 271 -56
rect 271 -57 272 -56
rect 272 -57 273 -56
rect 273 -57 274 -56
rect 274 -57 275 -56
rect 275 -57 276 -56
rect 276 -57 277 -56
rect 277 -57 278 -56
rect 278 -57 279 -56
rect 279 -57 280 -56
rect 280 -57 281 -56
rect 281 -57 282 -56
rect 282 -57 283 -56
rect 283 -57 284 -56
rect 284 -57 285 -56
rect 285 -57 286 -56
rect 286 -57 287 -56
rect 287 -57 288 -56
rect 288 -57 289 -56
rect 289 -57 290 -56
rect 290 -57 291 -56
rect 291 -57 292 -56
rect 292 -57 293 -56
rect 293 -57 294 -56
rect 294 -57 295 -56
rect 295 -57 296 -56
rect 296 -57 297 -56
rect 297 -57 298 -56
rect 298 -57 299 -56
rect 299 -57 300 -56
rect 300 -57 301 -56
rect 301 -57 302 -56
rect 302 -57 303 -56
rect 303 -57 304 -56
rect 304 -57 305 -56
rect 305 -57 306 -56
rect 306 -57 307 -56
rect 307 -57 308 -56
rect 308 -57 309 -56
rect 309 -57 310 -56
rect 310 -57 311 -56
rect 311 -57 312 -56
rect 312 -57 313 -56
rect 313 -57 314 -56
rect 314 -57 315 -56
rect 315 -57 316 -56
rect 316 -57 317 -56
rect 317 -57 318 -56
rect 318 -57 319 -56
rect 319 -57 320 -56
rect 320 -57 321 -56
rect 321 -57 322 -56
rect 322 -57 323 -56
rect 323 -57 324 -56
rect 324 -57 325 -56
rect 325 -57 326 -56
rect 326 -57 327 -56
rect 327 -57 328 -56
rect 328 -57 329 -56
rect 329 -57 330 -56
rect 330 -57 331 -56
rect 331 -57 332 -56
rect 332 -57 333 -56
rect 333 -57 334 -56
rect 334 -57 335 -56
rect 335 -57 336 -56
rect 336 -57 337 -56
rect 337 -57 338 -56
rect 338 -57 339 -56
rect 339 -57 340 -56
rect 340 -57 341 -56
rect 341 -57 342 -56
rect 342 -57 343 -56
rect 343 -57 344 -56
rect 344 -57 345 -56
rect 345 -57 346 -56
rect 346 -57 347 -56
rect 347 -57 348 -56
rect 348 -57 349 -56
rect 349 -57 350 -56
rect 350 -57 351 -56
rect 351 -57 352 -56
rect 352 -57 353 -56
rect 353 -57 354 -56
rect 354 -57 355 -56
rect 355 -57 356 -56
rect 356 -57 357 -56
rect 357 -57 358 -56
rect 358 -57 359 -56
rect 359 -57 360 -56
rect 360 -57 361 -56
rect 361 -57 362 -56
rect 362 -57 363 -56
rect 363 -57 364 -56
rect 364 -57 365 -56
rect 365 -57 366 -56
rect 366 -57 367 -56
rect 367 -57 368 -56
rect 368 -57 369 -56
rect 369 -57 370 -56
rect 370 -57 371 -56
rect 371 -57 372 -56
rect 372 -57 373 -56
rect 373 -57 374 -56
rect 374 -57 375 -56
rect 375 -57 376 -56
rect 376 -57 377 -56
rect 377 -57 378 -56
rect 378 -57 379 -56
rect 379 -57 380 -56
rect 380 -57 381 -56
rect 381 -57 382 -56
rect 382 -57 383 -56
rect 383 -57 384 -56
rect 384 -57 385 -56
rect 385 -57 386 -56
rect 386 -57 387 -56
rect 387 -57 388 -56
rect 388 -57 389 -56
rect 389 -57 390 -56
rect 390 -57 391 -56
rect 391 -57 392 -56
rect 392 -57 393 -56
rect 393 -57 394 -56
rect 394 -57 395 -56
rect 395 -57 396 -56
rect 396 -57 397 -56
rect 397 -57 398 -56
rect 398 -57 399 -56
rect 399 -57 400 -56
rect 400 -57 401 -56
rect 401 -57 402 -56
rect 402 -57 403 -56
rect 403 -57 404 -56
rect 404 -57 405 -56
rect 405 -57 406 -56
rect 406 -57 407 -56
rect 407 -57 408 -56
rect 408 -57 409 -56
rect 409 -57 410 -56
rect 410 -57 411 -56
rect 411 -57 412 -56
rect 412 -57 413 -56
rect 413 -57 414 -56
rect 414 -57 415 -56
rect 415 -57 416 -56
rect 416 -57 417 -56
rect 417 -57 418 -56
rect 418 -57 419 -56
rect 419 -57 420 -56
rect 420 -57 421 -56
rect 421 -57 422 -56
rect 422 -57 423 -56
rect 423 -57 424 -56
rect 424 -57 425 -56
rect 425 -57 426 -56
rect 426 -57 427 -56
rect 427 -57 428 -56
rect 428 -57 429 -56
rect 429 -57 430 -56
rect 430 -57 431 -56
rect 431 -57 432 -56
rect 432 -57 433 -56
rect 433 -57 434 -56
rect 434 -57 435 -56
rect 435 -57 436 -56
rect 436 -57 437 -56
rect 437 -57 438 -56
rect 438 -57 439 -56
rect 439 -57 440 -56
rect 440 -57 441 -56
rect 441 -57 442 -56
rect 442 -57 443 -56
rect 443 -57 444 -56
rect 444 -57 445 -56
rect 445 -57 446 -56
rect 446 -57 447 -56
rect 447 -57 448 -56
rect 448 -57 449 -56
rect 449 -57 450 -56
rect 450 -57 451 -56
rect 451 -57 452 -56
rect 452 -57 453 -56
rect 453 -57 454 -56
rect 454 -57 455 -56
rect 455 -57 456 -56
rect 456 -57 457 -56
rect 457 -57 458 -56
rect 458 -57 459 -56
rect 459 -57 460 -56
rect 460 -57 461 -56
rect 461 -57 462 -56
rect 462 -57 463 -56
rect 463 -57 464 -56
rect 464 -57 465 -56
rect 465 -57 466 -56
rect 466 -57 467 -56
rect 467 -57 468 -56
rect 468 -57 469 -56
rect 469 -57 470 -56
rect 470 -57 471 -56
rect 471 -57 472 -56
rect 472 -57 473 -56
rect 473 -57 474 -56
rect 474 -57 475 -56
rect 475 -57 476 -56
rect 476 -57 477 -56
rect 477 -57 478 -56
rect 478 -57 479 -56
rect 479 -57 480 -56
rect 2 -58 3 -57
rect 3 -58 4 -57
rect 4 -58 5 -57
rect 5 -58 6 -57
rect 6 -58 7 -57
rect 7 -58 8 -57
rect 8 -58 9 -57
rect 9 -58 10 -57
rect 10 -58 11 -57
rect 11 -58 12 -57
rect 12 -58 13 -57
rect 13 -58 14 -57
rect 14 -58 15 -57
rect 15 -58 16 -57
rect 16 -58 17 -57
rect 17 -58 18 -57
rect 18 -58 19 -57
rect 19 -58 20 -57
rect 20 -58 21 -57
rect 21 -58 22 -57
rect 22 -58 23 -57
rect 23 -58 24 -57
rect 24 -58 25 -57
rect 25 -58 26 -57
rect 26 -58 27 -57
rect 27 -58 28 -57
rect 37 -58 38 -57
rect 38 -58 39 -57
rect 39 -58 40 -57
rect 40 -58 41 -57
rect 41 -58 42 -57
rect 42 -58 43 -57
rect 43 -58 44 -57
rect 44 -58 45 -57
rect 45 -58 46 -57
rect 46 -58 47 -57
rect 47 -58 48 -57
rect 48 -58 49 -57
rect 49 -58 50 -57
rect 50 -58 51 -57
rect 51 -58 52 -57
rect 52 -58 53 -57
rect 53 -58 54 -57
rect 54 -58 55 -57
rect 55 -58 56 -57
rect 56 -58 57 -57
rect 57 -58 58 -57
rect 58 -58 59 -57
rect 59 -58 60 -57
rect 69 -58 70 -57
rect 70 -58 71 -57
rect 71 -58 72 -57
rect 72 -58 73 -57
rect 73 -58 74 -57
rect 74 -58 75 -57
rect 75 -58 76 -57
rect 76 -58 77 -57
rect 77 -58 78 -57
rect 78 -58 79 -57
rect 79 -58 80 -57
rect 80 -58 81 -57
rect 81 -58 82 -57
rect 82 -58 83 -57
rect 83 -58 84 -57
rect 84 -58 85 -57
rect 85 -58 86 -57
rect 86 -58 87 -57
rect 87 -58 88 -57
rect 88 -58 89 -57
rect 89 -58 90 -57
rect 90 -58 91 -57
rect 91 -58 92 -57
rect 101 -58 102 -57
rect 102 -58 103 -57
rect 103 -58 104 -57
rect 104 -58 105 -57
rect 105 -58 106 -57
rect 106 -58 107 -57
rect 107 -58 108 -57
rect 108 -58 109 -57
rect 109 -58 110 -57
rect 110 -58 111 -57
rect 111 -58 112 -57
rect 112 -58 113 -57
rect 113 -58 114 -57
rect 114 -58 115 -57
rect 115 -58 116 -57
rect 116 -58 117 -57
rect 117 -58 118 -57
rect 118 -58 119 -57
rect 119 -58 120 -57
rect 120 -58 121 -57
rect 121 -58 122 -57
rect 122 -58 123 -57
rect 123 -58 124 -57
rect 133 -58 134 -57
rect 134 -58 135 -57
rect 135 -58 136 -57
rect 136 -58 137 -57
rect 137 -58 138 -57
rect 138 -58 139 -57
rect 139 -58 140 -57
rect 140 -58 141 -57
rect 141 -58 142 -57
rect 142 -58 143 -57
rect 143 -58 144 -57
rect 144 -58 145 -57
rect 145 -58 146 -57
rect 146 -58 147 -57
rect 147 -58 148 -57
rect 148 -58 149 -57
rect 149 -58 150 -57
rect 150 -58 151 -57
rect 151 -58 152 -57
rect 152 -58 153 -57
rect 153 -58 154 -57
rect 154 -58 155 -57
rect 155 -58 156 -57
rect 165 -58 166 -57
rect 166 -58 167 -57
rect 167 -58 168 -57
rect 168 -58 169 -57
rect 169 -58 170 -57
rect 170 -58 171 -57
rect 171 -58 172 -57
rect 172 -58 173 -57
rect 173 -58 174 -57
rect 174 -58 175 -57
rect 175 -58 176 -57
rect 176 -58 177 -57
rect 177 -58 178 -57
rect 178 -58 179 -57
rect 179 -58 180 -57
rect 180 -58 181 -57
rect 181 -58 182 -57
rect 182 -58 183 -57
rect 183 -58 184 -57
rect 184 -58 185 -57
rect 185 -58 186 -57
rect 186 -58 187 -57
rect 187 -58 188 -57
rect 188 -58 189 -57
rect 189 -58 190 -57
rect 190 -58 191 -57
rect 191 -58 192 -57
rect 2 -59 3 -58
rect 3 -59 4 -58
rect 4 -59 5 -58
rect 5 -59 6 -58
rect 6 -59 7 -58
rect 7 -59 8 -58
rect 8 -59 9 -58
rect 9 -59 10 -58
rect 10 -59 11 -58
rect 11 -59 12 -58
rect 12 -59 13 -58
rect 13 -59 14 -58
rect 14 -59 15 -58
rect 15 -59 16 -58
rect 16 -59 17 -58
rect 17 -59 18 -58
rect 18 -59 19 -58
rect 19 -59 20 -58
rect 20 -59 21 -58
rect 21 -59 22 -58
rect 22 -59 23 -58
rect 23 -59 24 -58
rect 24 -59 25 -58
rect 25 -59 26 -58
rect 26 -59 27 -58
rect 27 -59 28 -58
rect 32 -59 33 -58
rect 33 -59 34 -58
rect 38 -59 39 -58
rect 39 -59 40 -58
rect 40 -59 41 -58
rect 41 -59 42 -58
rect 42 -59 43 -58
rect 43 -59 44 -58
rect 44 -59 45 -58
rect 45 -59 46 -58
rect 46 -59 47 -58
rect 47 -59 48 -58
rect 48 -59 49 -58
rect 49 -59 50 -58
rect 50 -59 51 -58
rect 51 -59 52 -58
rect 52 -59 53 -58
rect 53 -59 54 -58
rect 54 -59 55 -58
rect 55 -59 56 -58
rect 56 -59 57 -58
rect 57 -59 58 -58
rect 58 -59 59 -58
rect 59 -59 60 -58
rect 64 -59 65 -58
rect 65 -59 66 -58
rect 70 -59 71 -58
rect 71 -59 72 -58
rect 72 -59 73 -58
rect 73 -59 74 -58
rect 74 -59 75 -58
rect 75 -59 76 -58
rect 76 -59 77 -58
rect 77 -59 78 -58
rect 78 -59 79 -58
rect 79 -59 80 -58
rect 80 -59 81 -58
rect 81 -59 82 -58
rect 82 -59 83 -58
rect 83 -59 84 -58
rect 84 -59 85 -58
rect 85 -59 86 -58
rect 86 -59 87 -58
rect 87 -59 88 -58
rect 88 -59 89 -58
rect 89 -59 90 -58
rect 90 -59 91 -58
rect 91 -59 92 -58
rect 96 -59 97 -58
rect 97 -59 98 -58
rect 102 -59 103 -58
rect 103 -59 104 -58
rect 104 -59 105 -58
rect 105 -59 106 -58
rect 106 -59 107 -58
rect 107 -59 108 -58
rect 108 -59 109 -58
rect 109 -59 110 -58
rect 110 -59 111 -58
rect 111 -59 112 -58
rect 112 -59 113 -58
rect 113 -59 114 -58
rect 114 -59 115 -58
rect 115 -59 116 -58
rect 116 -59 117 -58
rect 117 -59 118 -58
rect 118 -59 119 -58
rect 119 -59 120 -58
rect 120 -59 121 -58
rect 121 -59 122 -58
rect 122 -59 123 -58
rect 123 -59 124 -58
rect 128 -59 129 -58
rect 129 -59 130 -58
rect 134 -59 135 -58
rect 135 -59 136 -58
rect 136 -59 137 -58
rect 137 -59 138 -58
rect 138 -59 139 -58
rect 139 -59 140 -58
rect 140 -59 141 -58
rect 141 -59 142 -58
rect 142 -59 143 -58
rect 143 -59 144 -58
rect 144 -59 145 -58
rect 145 -59 146 -58
rect 146 -59 147 -58
rect 147 -59 148 -58
rect 148 -59 149 -58
rect 149 -59 150 -58
rect 150 -59 151 -58
rect 151 -59 152 -58
rect 152 -59 153 -58
rect 153 -59 154 -58
rect 154 -59 155 -58
rect 155 -59 156 -58
rect 160 -59 161 -58
rect 161 -59 162 -58
rect 166 -59 167 -58
rect 167 -59 168 -58
rect 168 -59 169 -58
rect 169 -59 170 -58
rect 170 -59 171 -58
rect 171 -59 172 -58
rect 172 -59 173 -58
rect 173 -59 174 -58
rect 174 -59 175 -58
rect 175 -59 176 -58
rect 176 -59 177 -58
rect 177 -59 178 -58
rect 178 -59 179 -58
rect 179 -59 180 -58
rect 180 -59 181 -58
rect 181 -59 182 -58
rect 182 -59 183 -58
rect 183 -59 184 -58
rect 184 -59 185 -58
rect 185 -59 186 -58
rect 186 -59 187 -58
rect 187 -59 188 -58
rect 188 -59 189 -58
rect 189 -59 190 -58
rect 190 -59 191 -58
rect 191 -59 192 -58
rect 2 -60 3 -59
rect 3 -60 4 -59
rect 4 -60 5 -59
rect 5 -60 6 -59
rect 6 -60 7 -59
rect 7 -60 8 -59
rect 8 -60 9 -59
rect 9 -60 10 -59
rect 10 -60 11 -59
rect 11 -60 12 -59
rect 12 -60 13 -59
rect 13 -60 14 -59
rect 14 -60 15 -59
rect 15 -60 16 -59
rect 18 -60 19 -59
rect 19 -60 20 -59
rect 20 -60 21 -59
rect 21 -60 22 -59
rect 22 -60 23 -59
rect 23 -60 24 -59
rect 24 -60 25 -59
rect 25 -60 26 -59
rect 26 -60 27 -59
rect 27 -60 28 -59
rect 31 -60 32 -59
rect 32 -60 33 -59
rect 33 -60 34 -59
rect 34 -60 35 -59
rect 38 -60 39 -59
rect 39 -60 40 -59
rect 40 -60 41 -59
rect 41 -60 42 -59
rect 42 -60 43 -59
rect 43 -60 44 -59
rect 44 -60 45 -59
rect 45 -60 46 -59
rect 46 -60 47 -59
rect 47 -60 48 -59
rect 50 -60 51 -59
rect 51 -60 52 -59
rect 52 -60 53 -59
rect 53 -60 54 -59
rect 54 -60 55 -59
rect 55 -60 56 -59
rect 56 -60 57 -59
rect 57 -60 58 -59
rect 58 -60 59 -59
rect 59 -60 60 -59
rect 63 -60 64 -59
rect 64 -60 65 -59
rect 65 -60 66 -59
rect 66 -60 67 -59
rect 70 -60 71 -59
rect 71 -60 72 -59
rect 72 -60 73 -59
rect 73 -60 74 -59
rect 74 -60 75 -59
rect 75 -60 76 -59
rect 76 -60 77 -59
rect 77 -60 78 -59
rect 78 -60 79 -59
rect 79 -60 80 -59
rect 82 -60 83 -59
rect 83 -60 84 -59
rect 84 -60 85 -59
rect 85 -60 86 -59
rect 86 -60 87 -59
rect 87 -60 88 -59
rect 88 -60 89 -59
rect 89 -60 90 -59
rect 90 -60 91 -59
rect 91 -60 92 -59
rect 95 -60 96 -59
rect 96 -60 97 -59
rect 97 -60 98 -59
rect 98 -60 99 -59
rect 102 -60 103 -59
rect 103 -60 104 -59
rect 104 -60 105 -59
rect 105 -60 106 -59
rect 106 -60 107 -59
rect 107 -60 108 -59
rect 108 -60 109 -59
rect 109 -60 110 -59
rect 110 -60 111 -59
rect 111 -60 112 -59
rect 114 -60 115 -59
rect 115 -60 116 -59
rect 116 -60 117 -59
rect 117 -60 118 -59
rect 118 -60 119 -59
rect 119 -60 120 -59
rect 120 -60 121 -59
rect 121 -60 122 -59
rect 122 -60 123 -59
rect 123 -60 124 -59
rect 127 -60 128 -59
rect 128 -60 129 -59
rect 129 -60 130 -59
rect 130 -60 131 -59
rect 134 -60 135 -59
rect 135 -60 136 -59
rect 136 -60 137 -59
rect 137 -60 138 -59
rect 138 -60 139 -59
rect 139 -60 140 -59
rect 140 -60 141 -59
rect 141 -60 142 -59
rect 142 -60 143 -59
rect 143 -60 144 -59
rect 146 -60 147 -59
rect 147 -60 148 -59
rect 148 -60 149 -59
rect 149 -60 150 -59
rect 150 -60 151 -59
rect 151 -60 152 -59
rect 152 -60 153 -59
rect 153 -60 154 -59
rect 154 -60 155 -59
rect 155 -60 156 -59
rect 159 -60 160 -59
rect 160 -60 161 -59
rect 161 -60 162 -59
rect 162 -60 163 -59
rect 166 -60 167 -59
rect 167 -60 168 -59
rect 168 -60 169 -59
rect 169 -60 170 -59
rect 170 -60 171 -59
rect 171 -60 172 -59
rect 172 -60 173 -59
rect 173 -60 174 -59
rect 174 -60 175 -59
rect 175 -60 176 -59
rect 178 -60 179 -59
rect 179 -60 180 -59
rect 180 -60 181 -59
rect 181 -60 182 -59
rect 182 -60 183 -59
rect 183 -60 184 -59
rect 184 -60 185 -59
rect 185 -60 186 -59
rect 186 -60 187 -59
rect 187 -60 188 -59
rect 188 -60 189 -59
rect 189 -60 190 -59
rect 190 -60 191 -59
rect 191 -60 192 -59
rect 2 -61 3 -60
rect 3 -61 4 -60
rect 4 -61 5 -60
rect 5 -61 6 -60
rect 6 -61 7 -60
rect 7 -61 8 -60
rect 8 -61 9 -60
rect 9 -61 10 -60
rect 10 -61 11 -60
rect 11 -61 12 -60
rect 12 -61 13 -60
rect 13 -61 14 -60
rect 14 -61 15 -60
rect 18 -61 19 -60
rect 19 -61 20 -60
rect 20 -61 21 -60
rect 21 -61 22 -60
rect 22 -61 23 -60
rect 23 -61 24 -60
rect 24 -61 25 -60
rect 25 -61 26 -60
rect 26 -61 27 -60
rect 27 -61 28 -60
rect 28 -61 29 -60
rect 29 -61 30 -60
rect 30 -61 31 -60
rect 31 -61 32 -60
rect 32 -61 33 -60
rect 33 -61 34 -60
rect 34 -61 35 -60
rect 35 -61 36 -60
rect 36 -61 37 -60
rect 37 -61 38 -60
rect 38 -61 39 -60
rect 39 -61 40 -60
rect 40 -61 41 -60
rect 41 -61 42 -60
rect 42 -61 43 -60
rect 43 -61 44 -60
rect 44 -61 45 -60
rect 45 -61 46 -60
rect 46 -61 47 -60
rect 50 -61 51 -60
rect 51 -61 52 -60
rect 52 -61 53 -60
rect 53 -61 54 -60
rect 54 -61 55 -60
rect 55 -61 56 -60
rect 56 -61 57 -60
rect 57 -61 58 -60
rect 58 -61 59 -60
rect 59 -61 60 -60
rect 60 -61 61 -60
rect 61 -61 62 -60
rect 62 -61 63 -60
rect 63 -61 64 -60
rect 64 -61 65 -60
rect 65 -61 66 -60
rect 66 -61 67 -60
rect 67 -61 68 -60
rect 68 -61 69 -60
rect 69 -61 70 -60
rect 70 -61 71 -60
rect 71 -61 72 -60
rect 72 -61 73 -60
rect 73 -61 74 -60
rect 74 -61 75 -60
rect 75 -61 76 -60
rect 76 -61 77 -60
rect 77 -61 78 -60
rect 78 -61 79 -60
rect 82 -61 83 -60
rect 83 -61 84 -60
rect 84 -61 85 -60
rect 85 -61 86 -60
rect 86 -61 87 -60
rect 87 -61 88 -60
rect 88 -61 89 -60
rect 89 -61 90 -60
rect 90 -61 91 -60
rect 91 -61 92 -60
rect 92 -61 93 -60
rect 93 -61 94 -60
rect 94 -61 95 -60
rect 95 -61 96 -60
rect 96 -61 97 -60
rect 97 -61 98 -60
rect 98 -61 99 -60
rect 99 -61 100 -60
rect 100 -61 101 -60
rect 101 -61 102 -60
rect 102 -61 103 -60
rect 103 -61 104 -60
rect 104 -61 105 -60
rect 105 -61 106 -60
rect 106 -61 107 -60
rect 107 -61 108 -60
rect 108 -61 109 -60
rect 109 -61 110 -60
rect 110 -61 111 -60
rect 114 -61 115 -60
rect 115 -61 116 -60
rect 116 -61 117 -60
rect 117 -61 118 -60
rect 118 -61 119 -60
rect 119 -61 120 -60
rect 120 -61 121 -60
rect 121 -61 122 -60
rect 122 -61 123 -60
rect 123 -61 124 -60
rect 124 -61 125 -60
rect 125 -61 126 -60
rect 126 -61 127 -60
rect 127 -61 128 -60
rect 128 -61 129 -60
rect 129 -61 130 -60
rect 130 -61 131 -60
rect 131 -61 132 -60
rect 132 -61 133 -60
rect 133 -61 134 -60
rect 134 -61 135 -60
rect 135 -61 136 -60
rect 136 -61 137 -60
rect 137 -61 138 -60
rect 138 -61 139 -60
rect 139 -61 140 -60
rect 140 -61 141 -60
rect 141 -61 142 -60
rect 142 -61 143 -60
rect 146 -61 147 -60
rect 147 -61 148 -60
rect 148 -61 149 -60
rect 149 -61 150 -60
rect 150 -61 151 -60
rect 151 -61 152 -60
rect 152 -61 153 -60
rect 153 -61 154 -60
rect 154 -61 155 -60
rect 155 -61 156 -60
rect 156 -61 157 -60
rect 157 -61 158 -60
rect 158 -61 159 -60
rect 159 -61 160 -60
rect 160 -61 161 -60
rect 161 -61 162 -60
rect 162 -61 163 -60
rect 163 -61 164 -60
rect 164 -61 165 -60
rect 165 -61 166 -60
rect 166 -61 167 -60
rect 167 -61 168 -60
rect 168 -61 169 -60
rect 169 -61 170 -60
rect 170 -61 171 -60
rect 171 -61 172 -60
rect 172 -61 173 -60
rect 173 -61 174 -60
rect 174 -61 175 -60
rect 178 -61 179 -60
rect 179 -61 180 -60
rect 180 -61 181 -60
rect 181 -61 182 -60
rect 182 -61 183 -60
rect 183 -61 184 -60
rect 184 -61 185 -60
rect 185 -61 186 -60
rect 186 -61 187 -60
rect 187 -61 188 -60
rect 188 -61 189 -60
rect 189 -61 190 -60
rect 190 -61 191 -60
rect 191 -61 192 -60
rect 2 -62 3 -61
rect 3 -62 4 -61
rect 4 -62 5 -61
rect 5 -62 6 -61
rect 6 -62 7 -61
rect 7 -62 8 -61
rect 8 -62 9 -61
rect 9 -62 10 -61
rect 10 -62 11 -61
rect 11 -62 12 -61
rect 12 -62 13 -61
rect 13 -62 14 -61
rect 14 -62 15 -61
rect 19 -62 20 -61
rect 20 -62 21 -61
rect 21 -62 22 -61
rect 22 -62 23 -61
rect 23 -62 24 -61
rect 24 -62 25 -61
rect 25 -62 26 -61
rect 26 -62 27 -61
rect 27 -62 28 -61
rect 28 -62 29 -61
rect 29 -62 30 -61
rect 30 -62 31 -61
rect 31 -62 32 -61
rect 32 -62 33 -61
rect 33 -62 34 -61
rect 34 -62 35 -61
rect 35 -62 36 -61
rect 36 -62 37 -61
rect 37 -62 38 -61
rect 38 -62 39 -61
rect 39 -62 40 -61
rect 40 -62 41 -61
rect 41 -62 42 -61
rect 42 -62 43 -61
rect 43 -62 44 -61
rect 44 -62 45 -61
rect 45 -62 46 -61
rect 46 -62 47 -61
rect 51 -62 52 -61
rect 52 -62 53 -61
rect 53 -62 54 -61
rect 54 -62 55 -61
rect 55 -62 56 -61
rect 56 -62 57 -61
rect 57 -62 58 -61
rect 58 -62 59 -61
rect 59 -62 60 -61
rect 60 -62 61 -61
rect 61 -62 62 -61
rect 62 -62 63 -61
rect 63 -62 64 -61
rect 64 -62 65 -61
rect 65 -62 66 -61
rect 66 -62 67 -61
rect 67 -62 68 -61
rect 68 -62 69 -61
rect 69 -62 70 -61
rect 70 -62 71 -61
rect 71 -62 72 -61
rect 72 -62 73 -61
rect 73 -62 74 -61
rect 74 -62 75 -61
rect 75 -62 76 -61
rect 76 -62 77 -61
rect 77 -62 78 -61
rect 78 -62 79 -61
rect 83 -62 84 -61
rect 84 -62 85 -61
rect 85 -62 86 -61
rect 86 -62 87 -61
rect 87 -62 88 -61
rect 88 -62 89 -61
rect 89 -62 90 -61
rect 90 -62 91 -61
rect 91 -62 92 -61
rect 92 -62 93 -61
rect 93 -62 94 -61
rect 94 -62 95 -61
rect 95 -62 96 -61
rect 96 -62 97 -61
rect 97 -62 98 -61
rect 98 -62 99 -61
rect 99 -62 100 -61
rect 100 -62 101 -61
rect 101 -62 102 -61
rect 102 -62 103 -61
rect 103 -62 104 -61
rect 104 -62 105 -61
rect 105 -62 106 -61
rect 106 -62 107 -61
rect 107 -62 108 -61
rect 108 -62 109 -61
rect 109 -62 110 -61
rect 110 -62 111 -61
rect 115 -62 116 -61
rect 116 -62 117 -61
rect 117 -62 118 -61
rect 118 -62 119 -61
rect 119 -62 120 -61
rect 120 -62 121 -61
rect 121 -62 122 -61
rect 122 -62 123 -61
rect 123 -62 124 -61
rect 124 -62 125 -61
rect 125 -62 126 -61
rect 126 -62 127 -61
rect 127 -62 128 -61
rect 128 -62 129 -61
rect 129 -62 130 -61
rect 130 -62 131 -61
rect 131 -62 132 -61
rect 132 -62 133 -61
rect 133 -62 134 -61
rect 134 -62 135 -61
rect 135 -62 136 -61
rect 136 -62 137 -61
rect 137 -62 138 -61
rect 138 -62 139 -61
rect 139 -62 140 -61
rect 140 -62 141 -61
rect 141 -62 142 -61
rect 142 -62 143 -61
rect 147 -62 148 -61
rect 148 -62 149 -61
rect 149 -62 150 -61
rect 150 -62 151 -61
rect 151 -62 152 -61
rect 152 -62 153 -61
rect 153 -62 154 -61
rect 154 -62 155 -61
rect 155 -62 156 -61
rect 156 -62 157 -61
rect 157 -62 158 -61
rect 158 -62 159 -61
rect 159 -62 160 -61
rect 160 -62 161 -61
rect 161 -62 162 -61
rect 162 -62 163 -61
rect 163 -62 164 -61
rect 164 -62 165 -61
rect 165 -62 166 -61
rect 166 -62 167 -61
rect 167 -62 168 -61
rect 168 -62 169 -61
rect 169 -62 170 -61
rect 170 -62 171 -61
rect 171 -62 172 -61
rect 172 -62 173 -61
rect 173 -62 174 -61
rect 174 -62 175 -61
rect 179 -62 180 -61
rect 180 -62 181 -61
rect 181 -62 182 -61
rect 182 -62 183 -61
rect 183 -62 184 -61
rect 184 -62 185 -61
rect 185 -62 186 -61
rect 186 -62 187 -61
rect 187 -62 188 -61
rect 188 -62 189 -61
rect 189 -62 190 -61
rect 190 -62 191 -61
rect 191 -62 192 -61
rect 2 -63 3 -62
rect 3 -63 4 -62
rect 4 -63 5 -62
rect 5 -63 6 -62
rect 6 -63 7 -62
rect 7 -63 8 -62
rect 8 -63 9 -62
rect 9 -63 10 -62
rect 10 -63 11 -62
rect 11 -63 12 -62
rect 12 -63 13 -62
rect 13 -63 14 -62
rect 14 -63 15 -62
rect 19 -63 20 -62
rect 20 -63 21 -62
rect 21 -63 22 -62
rect 22 -63 23 -62
rect 23 -63 24 -62
rect 24 -63 25 -62
rect 25 -63 26 -62
rect 26 -63 27 -62
rect 27 -63 28 -62
rect 28 -63 29 -62
rect 29 -63 30 -62
rect 30 -63 31 -62
rect 31 -63 32 -62
rect 32 -63 33 -62
rect 33 -63 34 -62
rect 34 -63 35 -62
rect 35 -63 36 -62
rect 36 -63 37 -62
rect 37 -63 38 -62
rect 38 -63 39 -62
rect 39 -63 40 -62
rect 40 -63 41 -62
rect 41 -63 42 -62
rect 42 -63 43 -62
rect 43 -63 44 -62
rect 44 -63 45 -62
rect 45 -63 46 -62
rect 46 -63 47 -62
rect 51 -63 52 -62
rect 52 -63 53 -62
rect 53 -63 54 -62
rect 54 -63 55 -62
rect 55 -63 56 -62
rect 56 -63 57 -62
rect 57 -63 58 -62
rect 58 -63 59 -62
rect 59 -63 60 -62
rect 60 -63 61 -62
rect 61 -63 62 -62
rect 62 -63 63 -62
rect 63 -63 64 -62
rect 64 -63 65 -62
rect 65 -63 66 -62
rect 66 -63 67 -62
rect 67 -63 68 -62
rect 68 -63 69 -62
rect 69 -63 70 -62
rect 70 -63 71 -62
rect 71 -63 72 -62
rect 72 -63 73 -62
rect 73 -63 74 -62
rect 74 -63 75 -62
rect 75 -63 76 -62
rect 76 -63 77 -62
rect 77 -63 78 -62
rect 78 -63 79 -62
rect 83 -63 84 -62
rect 84 -63 85 -62
rect 85 -63 86 -62
rect 86 -63 87 -62
rect 87 -63 88 -62
rect 88 -63 89 -62
rect 89 -63 90 -62
rect 90 -63 91 -62
rect 91 -63 92 -62
rect 92 -63 93 -62
rect 93 -63 94 -62
rect 94 -63 95 -62
rect 95 -63 96 -62
rect 96 -63 97 -62
rect 97 -63 98 -62
rect 98 -63 99 -62
rect 99 -63 100 -62
rect 100 -63 101 -62
rect 101 -63 102 -62
rect 102 -63 103 -62
rect 103 -63 104 -62
rect 104 -63 105 -62
rect 105 -63 106 -62
rect 106 -63 107 -62
rect 107 -63 108 -62
rect 108 -63 109 -62
rect 109 -63 110 -62
rect 110 -63 111 -62
rect 115 -63 116 -62
rect 116 -63 117 -62
rect 117 -63 118 -62
rect 118 -63 119 -62
rect 119 -63 120 -62
rect 120 -63 121 -62
rect 121 -63 122 -62
rect 122 -63 123 -62
rect 123 -63 124 -62
rect 124 -63 125 -62
rect 125 -63 126 -62
rect 126 -63 127 -62
rect 127 -63 128 -62
rect 128 -63 129 -62
rect 129 -63 130 -62
rect 130 -63 131 -62
rect 131 -63 132 -62
rect 132 -63 133 -62
rect 133 -63 134 -62
rect 134 -63 135 -62
rect 135 -63 136 -62
rect 136 -63 137 -62
rect 137 -63 138 -62
rect 138 -63 139 -62
rect 139 -63 140 -62
rect 140 -63 141 -62
rect 141 -63 142 -62
rect 142 -63 143 -62
rect 147 -63 148 -62
rect 148 -63 149 -62
rect 149 -63 150 -62
rect 150 -63 151 -62
rect 151 -63 152 -62
rect 152 -63 153 -62
rect 153 -63 154 -62
rect 154 -63 155 -62
rect 155 -63 156 -62
rect 156 -63 157 -62
rect 157 -63 158 -62
rect 158 -63 159 -62
rect 159 -63 160 -62
rect 160 -63 161 -62
rect 161 -63 162 -62
rect 162 -63 163 -62
rect 163 -63 164 -62
rect 164 -63 165 -62
rect 165 -63 166 -62
rect 166 -63 167 -62
rect 167 -63 168 -62
rect 168 -63 169 -62
rect 169 -63 170 -62
rect 170 -63 171 -62
rect 171 -63 172 -62
rect 172 -63 173 -62
rect 173 -63 174 -62
rect 174 -63 175 -62
rect 179 -63 180 -62
rect 180 -63 181 -62
rect 181 -63 182 -62
rect 182 -63 183 -62
rect 183 -63 184 -62
rect 184 -63 185 -62
rect 185 -63 186 -62
rect 186 -63 187 -62
rect 187 -63 188 -62
rect 188 -63 189 -62
rect 189 -63 190 -62
rect 190 -63 191 -62
rect 191 -63 192 -62
rect 2 -64 3 -63
rect 3 -64 4 -63
rect 4 -64 5 -63
rect 5 -64 6 -63
rect 6 -64 7 -63
rect 7 -64 8 -63
rect 8 -64 9 -63
rect 9 -64 10 -63
rect 10 -64 11 -63
rect 11 -64 12 -63
rect 12 -64 13 -63
rect 13 -64 14 -63
rect 19 -64 20 -63
rect 20 -64 21 -63
rect 21 -64 22 -63
rect 22 -64 23 -63
rect 23 -64 24 -63
rect 24 -64 25 -63
rect 25 -64 26 -63
rect 26 -64 27 -63
rect 27 -64 28 -63
rect 28 -64 29 -63
rect 29 -64 30 -63
rect 30 -64 31 -63
rect 31 -64 32 -63
rect 32 -64 33 -63
rect 33 -64 34 -63
rect 34 -64 35 -63
rect 35 -64 36 -63
rect 36 -64 37 -63
rect 37 -64 38 -63
rect 38 -64 39 -63
rect 39 -64 40 -63
rect 40 -64 41 -63
rect 41 -64 42 -63
rect 42 -64 43 -63
rect 43 -64 44 -63
rect 44 -64 45 -63
rect 45 -64 46 -63
rect 51 -64 52 -63
rect 52 -64 53 -63
rect 53 -64 54 -63
rect 54 -64 55 -63
rect 55 -64 56 -63
rect 56 -64 57 -63
rect 57 -64 58 -63
rect 58 -64 59 -63
rect 59 -64 60 -63
rect 60 -64 61 -63
rect 61 -64 62 -63
rect 62 -64 63 -63
rect 63 -64 64 -63
rect 64 -64 65 -63
rect 65 -64 66 -63
rect 66 -64 67 -63
rect 67 -64 68 -63
rect 68 -64 69 -63
rect 69 -64 70 -63
rect 70 -64 71 -63
rect 71 -64 72 -63
rect 72 -64 73 -63
rect 73 -64 74 -63
rect 74 -64 75 -63
rect 75 -64 76 -63
rect 76 -64 77 -63
rect 77 -64 78 -63
rect 83 -64 84 -63
rect 84 -64 85 -63
rect 85 -64 86 -63
rect 86 -64 87 -63
rect 87 -64 88 -63
rect 88 -64 89 -63
rect 89 -64 90 -63
rect 90 -64 91 -63
rect 91 -64 92 -63
rect 92 -64 93 -63
rect 93 -64 94 -63
rect 94 -64 95 -63
rect 95 -64 96 -63
rect 96 -64 97 -63
rect 97 -64 98 -63
rect 98 -64 99 -63
rect 99 -64 100 -63
rect 100 -64 101 -63
rect 101 -64 102 -63
rect 102 -64 103 -63
rect 103 -64 104 -63
rect 104 -64 105 -63
rect 105 -64 106 -63
rect 106 -64 107 -63
rect 107 -64 108 -63
rect 108 -64 109 -63
rect 109 -64 110 -63
rect 115 -64 116 -63
rect 116 -64 117 -63
rect 117 -64 118 -63
rect 118 -64 119 -63
rect 119 -64 120 -63
rect 120 -64 121 -63
rect 121 -64 122 -63
rect 122 -64 123 -63
rect 123 -64 124 -63
rect 124 -64 125 -63
rect 125 -64 126 -63
rect 126 -64 127 -63
rect 127 -64 128 -63
rect 128 -64 129 -63
rect 129 -64 130 -63
rect 130 -64 131 -63
rect 131 -64 132 -63
rect 132 -64 133 -63
rect 133 -64 134 -63
rect 134 -64 135 -63
rect 135 -64 136 -63
rect 136 -64 137 -63
rect 137 -64 138 -63
rect 138 -64 139 -63
rect 139 -64 140 -63
rect 140 -64 141 -63
rect 141 -64 142 -63
rect 147 -64 148 -63
rect 148 -64 149 -63
rect 149 -64 150 -63
rect 150 -64 151 -63
rect 151 -64 152 -63
rect 152 -64 153 -63
rect 153 -64 154 -63
rect 154 -64 155 -63
rect 155 -64 156 -63
rect 156 -64 157 -63
rect 157 -64 158 -63
rect 158 -64 159 -63
rect 159 -64 160 -63
rect 160 -64 161 -63
rect 161 -64 162 -63
rect 162 -64 163 -63
rect 163 -64 164 -63
rect 164 -64 165 -63
rect 165 -64 166 -63
rect 166 -64 167 -63
rect 167 -64 168 -63
rect 168 -64 169 -63
rect 169 -64 170 -63
rect 170 -64 171 -63
rect 171 -64 172 -63
rect 172 -64 173 -63
rect 173 -64 174 -63
rect 179 -64 180 -63
rect 180 -64 181 -63
rect 181 -64 182 -63
rect 182 -64 183 -63
rect 183 -64 184 -63
rect 184 -64 185 -63
rect 185 -64 186 -63
rect 186 -64 187 -63
rect 187 -64 188 -63
rect 188 -64 189 -63
rect 189 -64 190 -63
rect 190 -64 191 -63
rect 191 -64 192 -63
rect 2 -65 3 -64
rect 3 -65 4 -64
rect 4 -65 5 -64
rect 5 -65 6 -64
rect 6 -65 7 -64
rect 7 -65 8 -64
rect 8 -65 9 -64
rect 25 -65 26 -64
rect 26 -65 27 -64
rect 27 -65 28 -64
rect 28 -65 29 -64
rect 29 -65 30 -64
rect 30 -65 31 -64
rect 31 -65 32 -64
rect 32 -65 33 -64
rect 33 -65 34 -64
rect 34 -65 35 -64
rect 35 -65 36 -64
rect 36 -65 37 -64
rect 37 -65 38 -64
rect 38 -65 39 -64
rect 39 -65 40 -64
rect 40 -65 41 -64
rect 57 -65 58 -64
rect 58 -65 59 -64
rect 59 -65 60 -64
rect 60 -65 61 -64
rect 61 -65 62 -64
rect 62 -65 63 -64
rect 63 -65 64 -64
rect 64 -65 65 -64
rect 65 -65 66 -64
rect 66 -65 67 -64
rect 67 -65 68 -64
rect 68 -65 69 -64
rect 69 -65 70 -64
rect 70 -65 71 -64
rect 71 -65 72 -64
rect 72 -65 73 -64
rect 89 -65 90 -64
rect 90 -65 91 -64
rect 91 -65 92 -64
rect 92 -65 93 -64
rect 93 -65 94 -64
rect 94 -65 95 -64
rect 95 -65 96 -64
rect 96 -65 97 -64
rect 97 -65 98 -64
rect 98 -65 99 -64
rect 99 -65 100 -64
rect 100 -65 101 -64
rect 101 -65 102 -64
rect 102 -65 103 -64
rect 103 -65 104 -64
rect 104 -65 105 -64
rect 121 -65 122 -64
rect 122 -65 123 -64
rect 123 -65 124 -64
rect 124 -65 125 -64
rect 125 -65 126 -64
rect 126 -65 127 -64
rect 127 -65 128 -64
rect 128 -65 129 -64
rect 129 -65 130 -64
rect 130 -65 131 -64
rect 131 -65 132 -64
rect 132 -65 133 -64
rect 133 -65 134 -64
rect 134 -65 135 -64
rect 135 -65 136 -64
rect 136 -65 137 -64
rect 153 -65 154 -64
rect 154 -65 155 -64
rect 155 -65 156 -64
rect 156 -65 157 -64
rect 157 -65 158 -64
rect 158 -65 159 -64
rect 159 -65 160 -64
rect 160 -65 161 -64
rect 161 -65 162 -64
rect 162 -65 163 -64
rect 163 -65 164 -64
rect 164 -65 165 -64
rect 165 -65 166 -64
rect 166 -65 167 -64
rect 167 -65 168 -64
rect 168 -65 169 -64
rect 185 -65 186 -64
rect 186 -65 187 -64
rect 187 -65 188 -64
rect 188 -65 189 -64
rect 189 -65 190 -64
rect 190 -65 191 -64
rect 191 -65 192 -64
rect 2 -66 3 -65
rect 3 -66 4 -65
rect 4 -66 5 -65
rect 5 -66 6 -65
rect 6 -66 7 -65
rect 7 -66 8 -65
rect 8 -66 9 -65
rect 25 -66 26 -65
rect 26 -66 27 -65
rect 27 -66 28 -65
rect 28 -66 29 -65
rect 29 -66 30 -65
rect 30 -66 31 -65
rect 31 -66 32 -65
rect 32 -66 33 -65
rect 33 -66 34 -65
rect 34 -66 35 -65
rect 35 -66 36 -65
rect 36 -66 37 -65
rect 37 -66 38 -65
rect 38 -66 39 -65
rect 39 -66 40 -65
rect 40 -66 41 -65
rect 57 -66 58 -65
rect 58 -66 59 -65
rect 59 -66 60 -65
rect 60 -66 61 -65
rect 61 -66 62 -65
rect 62 -66 63 -65
rect 63 -66 64 -65
rect 64 -66 65 -65
rect 65 -66 66 -65
rect 66 -66 67 -65
rect 67 -66 68 -65
rect 68 -66 69 -65
rect 69 -66 70 -65
rect 70 -66 71 -65
rect 71 -66 72 -65
rect 72 -66 73 -65
rect 89 -66 90 -65
rect 90 -66 91 -65
rect 91 -66 92 -65
rect 92 -66 93 -65
rect 93 -66 94 -65
rect 94 -66 95 -65
rect 95 -66 96 -65
rect 96 -66 97 -65
rect 97 -66 98 -65
rect 98 -66 99 -65
rect 99 -66 100 -65
rect 100 -66 101 -65
rect 101 -66 102 -65
rect 102 -66 103 -65
rect 103 -66 104 -65
rect 104 -66 105 -65
rect 121 -66 122 -65
rect 122 -66 123 -65
rect 123 -66 124 -65
rect 124 -66 125 -65
rect 125 -66 126 -65
rect 126 -66 127 -65
rect 127 -66 128 -65
rect 128 -66 129 -65
rect 129 -66 130 -65
rect 130 -66 131 -65
rect 131 -66 132 -65
rect 132 -66 133 -65
rect 133 -66 134 -65
rect 134 -66 135 -65
rect 135 -66 136 -65
rect 136 -66 137 -65
rect 153 -66 154 -65
rect 154 -66 155 -65
rect 155 -66 156 -65
rect 156 -66 157 -65
rect 157 -66 158 -65
rect 158 -66 159 -65
rect 159 -66 160 -65
rect 160 -66 161 -65
rect 161 -66 162 -65
rect 162 -66 163 -65
rect 163 -66 164 -65
rect 164 -66 165 -65
rect 165 -66 166 -65
rect 166 -66 167 -65
rect 167 -66 168 -65
rect 168 -66 169 -65
rect 185 -66 186 -65
rect 186 -66 187 -65
rect 187 -66 188 -65
rect 188 -66 189 -65
rect 189 -66 190 -65
rect 190 -66 191 -65
rect 191 -66 192 -65
rect 2 -67 3 -66
rect 3 -67 4 -66
rect 4 -67 5 -66
rect 5 -67 6 -66
rect 6 -67 7 -66
rect 7 -67 8 -66
rect 8 -67 9 -66
rect 9 -67 10 -66
rect 23 -67 24 -66
rect 24 -67 25 -66
rect 25 -67 26 -66
rect 26 -67 27 -66
rect 27 -67 28 -66
rect 28 -67 29 -66
rect 29 -67 30 -66
rect 30 -67 31 -66
rect 31 -67 32 -66
rect 32 -67 33 -66
rect 33 -67 34 -66
rect 34 -67 35 -66
rect 35 -67 36 -66
rect 36 -67 37 -66
rect 37 -67 38 -66
rect 38 -67 39 -66
rect 39 -67 40 -66
rect 40 -67 41 -66
rect 41 -67 42 -66
rect 55 -67 56 -66
rect 56 -67 57 -66
rect 57 -67 58 -66
rect 58 -67 59 -66
rect 59 -67 60 -66
rect 60 -67 61 -66
rect 61 -67 62 -66
rect 62 -67 63 -66
rect 63 -67 64 -66
rect 64 -67 65 -66
rect 65 -67 66 -66
rect 66 -67 67 -66
rect 67 -67 68 -66
rect 68 -67 69 -66
rect 69 -67 70 -66
rect 70 -67 71 -66
rect 71 -67 72 -66
rect 72 -67 73 -66
rect 73 -67 74 -66
rect 87 -67 88 -66
rect 88 -67 89 -66
rect 89 -67 90 -66
rect 90 -67 91 -66
rect 91 -67 92 -66
rect 92 -67 93 -66
rect 93 -67 94 -66
rect 94 -67 95 -66
rect 95 -67 96 -66
rect 96 -67 97 -66
rect 97 -67 98 -66
rect 98 -67 99 -66
rect 99 -67 100 -66
rect 100 -67 101 -66
rect 101 -67 102 -66
rect 102 -67 103 -66
rect 103 -67 104 -66
rect 104 -67 105 -66
rect 105 -67 106 -66
rect 119 -67 120 -66
rect 120 -67 121 -66
rect 121 -67 122 -66
rect 122 -67 123 -66
rect 123 -67 124 -66
rect 124 -67 125 -66
rect 125 -67 126 -66
rect 126 -67 127 -66
rect 127 -67 128 -66
rect 128 -67 129 -66
rect 129 -67 130 -66
rect 130 -67 131 -66
rect 131 -67 132 -66
rect 132 -67 133 -66
rect 133 -67 134 -66
rect 134 -67 135 -66
rect 135 -67 136 -66
rect 136 -67 137 -66
rect 137 -67 138 -66
rect 151 -67 152 -66
rect 152 -67 153 -66
rect 153 -67 154 -66
rect 154 -67 155 -66
rect 155 -67 156 -66
rect 156 -67 157 -66
rect 157 -67 158 -66
rect 158 -67 159 -66
rect 159 -67 160 -66
rect 160 -67 161 -66
rect 161 -67 162 -66
rect 162 -67 163 -66
rect 163 -67 164 -66
rect 164 -67 165 -66
rect 165 -67 166 -66
rect 166 -67 167 -66
rect 167 -67 168 -66
rect 168 -67 169 -66
rect 169 -67 170 -66
rect 183 -67 184 -66
rect 184 -67 185 -66
rect 185 -67 186 -66
rect 186 -67 187 -66
rect 187 -67 188 -66
rect 188 -67 189 -66
rect 189 -67 190 -66
rect 190 -67 191 -66
rect 191 -67 192 -66
rect 2 -68 3 -67
rect 3 -68 4 -67
rect 4 -68 5 -67
rect 5 -68 6 -67
rect 6 -68 7 -67
rect 7 -68 8 -67
rect 8 -68 9 -67
rect 9 -68 10 -67
rect 10 -68 11 -67
rect 22 -68 23 -67
rect 23 -68 24 -67
rect 24 -68 25 -67
rect 25 -68 26 -67
rect 26 -68 27 -67
rect 27 -68 28 -67
rect 28 -68 29 -67
rect 29 -68 30 -67
rect 30 -68 31 -67
rect 31 -68 32 -67
rect 32 -68 33 -67
rect 33 -68 34 -67
rect 34 -68 35 -67
rect 35 -68 36 -67
rect 36 -68 37 -67
rect 37 -68 38 -67
rect 38 -68 39 -67
rect 39 -68 40 -67
rect 40 -68 41 -67
rect 41 -68 42 -67
rect 42 -68 43 -67
rect 54 -68 55 -67
rect 55 -68 56 -67
rect 56 -68 57 -67
rect 57 -68 58 -67
rect 58 -68 59 -67
rect 59 -68 60 -67
rect 60 -68 61 -67
rect 61 -68 62 -67
rect 62 -68 63 -67
rect 63 -68 64 -67
rect 64 -68 65 -67
rect 65 -68 66 -67
rect 66 -68 67 -67
rect 67 -68 68 -67
rect 68 -68 69 -67
rect 69 -68 70 -67
rect 70 -68 71 -67
rect 71 -68 72 -67
rect 72 -68 73 -67
rect 73 -68 74 -67
rect 74 -68 75 -67
rect 86 -68 87 -67
rect 87 -68 88 -67
rect 88 -68 89 -67
rect 89 -68 90 -67
rect 90 -68 91 -67
rect 91 -68 92 -67
rect 92 -68 93 -67
rect 93 -68 94 -67
rect 94 -68 95 -67
rect 95 -68 96 -67
rect 96 -68 97 -67
rect 97 -68 98 -67
rect 98 -68 99 -67
rect 99 -68 100 -67
rect 100 -68 101 -67
rect 101 -68 102 -67
rect 102 -68 103 -67
rect 103 -68 104 -67
rect 104 -68 105 -67
rect 105 -68 106 -67
rect 106 -68 107 -67
rect 118 -68 119 -67
rect 119 -68 120 -67
rect 120 -68 121 -67
rect 121 -68 122 -67
rect 122 -68 123 -67
rect 123 -68 124 -67
rect 124 -68 125 -67
rect 125 -68 126 -67
rect 126 -68 127 -67
rect 127 -68 128 -67
rect 128 -68 129 -67
rect 129 -68 130 -67
rect 130 -68 131 -67
rect 131 -68 132 -67
rect 132 -68 133 -67
rect 133 -68 134 -67
rect 134 -68 135 -67
rect 135 -68 136 -67
rect 136 -68 137 -67
rect 137 -68 138 -67
rect 138 -68 139 -67
rect 150 -68 151 -67
rect 151 -68 152 -67
rect 152 -68 153 -67
rect 153 -68 154 -67
rect 154 -68 155 -67
rect 155 -68 156 -67
rect 156 -68 157 -67
rect 157 -68 158 -67
rect 158 -68 159 -67
rect 159 -68 160 -67
rect 160 -68 161 -67
rect 161 -68 162 -67
rect 162 -68 163 -67
rect 163 -68 164 -67
rect 164 -68 165 -67
rect 165 -68 166 -67
rect 166 -68 167 -67
rect 167 -68 168 -67
rect 168 -68 169 -67
rect 169 -68 170 -67
rect 170 -68 171 -67
rect 182 -68 183 -67
rect 183 -68 184 -67
rect 184 -68 185 -67
rect 185 -68 186 -67
rect 186 -68 187 -67
rect 187 -68 188 -67
rect 188 -68 189 -67
rect 189 -68 190 -67
rect 190 -68 191 -67
rect 191 -68 192 -67
rect 2 -69 3 -68
rect 3 -69 4 -68
rect 4 -69 5 -68
rect 5 -69 6 -68
rect 6 -69 7 -68
rect 7 -69 8 -68
rect 8 -69 9 -68
rect 9 -69 10 -68
rect 10 -69 11 -68
rect 11 -69 12 -68
rect 21 -69 22 -68
rect 22 -69 23 -68
rect 23 -69 24 -68
rect 24 -69 25 -68
rect 25 -69 26 -68
rect 26 -69 27 -68
rect 27 -69 28 -68
rect 28 -69 29 -68
rect 29 -69 30 -68
rect 30 -69 31 -68
rect 31 -69 32 -68
rect 32 -69 33 -68
rect 33 -69 34 -68
rect 34 -69 35 -68
rect 35 -69 36 -68
rect 36 -69 37 -68
rect 37 -69 38 -68
rect 38 -69 39 -68
rect 39 -69 40 -68
rect 40 -69 41 -68
rect 41 -69 42 -68
rect 42 -69 43 -68
rect 43 -69 44 -68
rect 53 -69 54 -68
rect 54 -69 55 -68
rect 55 -69 56 -68
rect 56 -69 57 -68
rect 57 -69 58 -68
rect 58 -69 59 -68
rect 59 -69 60 -68
rect 60 -69 61 -68
rect 61 -69 62 -68
rect 62 -69 63 -68
rect 63 -69 64 -68
rect 64 -69 65 -68
rect 65 -69 66 -68
rect 66 -69 67 -68
rect 67 -69 68 -68
rect 68 -69 69 -68
rect 69 -69 70 -68
rect 70 -69 71 -68
rect 71 -69 72 -68
rect 72 -69 73 -68
rect 73 -69 74 -68
rect 74 -69 75 -68
rect 75 -69 76 -68
rect 85 -69 86 -68
rect 86 -69 87 -68
rect 87 -69 88 -68
rect 88 -69 89 -68
rect 89 -69 90 -68
rect 90 -69 91 -68
rect 91 -69 92 -68
rect 92 -69 93 -68
rect 93 -69 94 -68
rect 94 -69 95 -68
rect 95 -69 96 -68
rect 96 -69 97 -68
rect 97 -69 98 -68
rect 98 -69 99 -68
rect 99 -69 100 -68
rect 100 -69 101 -68
rect 101 -69 102 -68
rect 102 -69 103 -68
rect 103 -69 104 -68
rect 104 -69 105 -68
rect 105 -69 106 -68
rect 106 -69 107 -68
rect 107 -69 108 -68
rect 117 -69 118 -68
rect 118 -69 119 -68
rect 119 -69 120 -68
rect 120 -69 121 -68
rect 121 -69 122 -68
rect 122 -69 123 -68
rect 123 -69 124 -68
rect 124 -69 125 -68
rect 125 -69 126 -68
rect 126 -69 127 -68
rect 127 -69 128 -68
rect 128 -69 129 -68
rect 129 -69 130 -68
rect 130 -69 131 -68
rect 131 -69 132 -68
rect 132 -69 133 -68
rect 133 -69 134 -68
rect 134 -69 135 -68
rect 135 -69 136 -68
rect 136 -69 137 -68
rect 137 -69 138 -68
rect 138 -69 139 -68
rect 139 -69 140 -68
rect 149 -69 150 -68
rect 150 -69 151 -68
rect 151 -69 152 -68
rect 152 -69 153 -68
rect 153 -69 154 -68
rect 154 -69 155 -68
rect 155 -69 156 -68
rect 156 -69 157 -68
rect 157 -69 158 -68
rect 158 -69 159 -68
rect 159 -69 160 -68
rect 160 -69 161 -68
rect 161 -69 162 -68
rect 162 -69 163 -68
rect 163 -69 164 -68
rect 164 -69 165 -68
rect 165 -69 166 -68
rect 166 -69 167 -68
rect 167 -69 168 -68
rect 168 -69 169 -68
rect 169 -69 170 -68
rect 170 -69 171 -68
rect 171 -69 172 -68
rect 181 -69 182 -68
rect 182 -69 183 -68
rect 183 -69 184 -68
rect 184 -69 185 -68
rect 185 -69 186 -68
rect 186 -69 187 -68
rect 187 -69 188 -68
rect 188 -69 189 -68
rect 189 -69 190 -68
rect 190 -69 191 -68
rect 191 -69 192 -68
rect 2 -70 3 -69
rect 3 -70 4 -69
rect 4 -70 5 -69
rect 5 -70 6 -69
rect 6 -70 7 -69
rect 7 -70 8 -69
rect 8 -70 9 -69
rect 9 -70 10 -69
rect 10 -70 11 -69
rect 11 -70 12 -69
rect 21 -70 22 -69
rect 22 -70 23 -69
rect 23 -70 24 -69
rect 24 -70 25 -69
rect 25 -70 26 -69
rect 26 -70 27 -69
rect 27 -70 28 -69
rect 28 -70 29 -69
rect 29 -70 30 -69
rect 30 -70 31 -69
rect 31 -70 32 -69
rect 32 -70 33 -69
rect 33 -70 34 -69
rect 34 -70 35 -69
rect 35 -70 36 -69
rect 36 -70 37 -69
rect 37 -70 38 -69
rect 38 -70 39 -69
rect 39 -70 40 -69
rect 40 -70 41 -69
rect 41 -70 42 -69
rect 42 -70 43 -69
rect 43 -70 44 -69
rect 53 -70 54 -69
rect 54 -70 55 -69
rect 55 -70 56 -69
rect 56 -70 57 -69
rect 57 -70 58 -69
rect 58 -70 59 -69
rect 59 -70 60 -69
rect 60 -70 61 -69
rect 61 -70 62 -69
rect 62 -70 63 -69
rect 63 -70 64 -69
rect 64 -70 65 -69
rect 65 -70 66 -69
rect 66 -70 67 -69
rect 67 -70 68 -69
rect 68 -70 69 -69
rect 69 -70 70 -69
rect 70 -70 71 -69
rect 71 -70 72 -69
rect 72 -70 73 -69
rect 73 -70 74 -69
rect 74 -70 75 -69
rect 75 -70 76 -69
rect 85 -70 86 -69
rect 86 -70 87 -69
rect 87 -70 88 -69
rect 88 -70 89 -69
rect 89 -70 90 -69
rect 90 -70 91 -69
rect 91 -70 92 -69
rect 92 -70 93 -69
rect 93 -70 94 -69
rect 94 -70 95 -69
rect 95 -70 96 -69
rect 96 -70 97 -69
rect 97 -70 98 -69
rect 98 -70 99 -69
rect 99 -70 100 -69
rect 100 -70 101 -69
rect 101 -70 102 -69
rect 102 -70 103 -69
rect 103 -70 104 -69
rect 104 -70 105 -69
rect 105 -70 106 -69
rect 106 -70 107 -69
rect 107 -70 108 -69
rect 117 -70 118 -69
rect 118 -70 119 -69
rect 119 -70 120 -69
rect 120 -70 121 -69
rect 121 -70 122 -69
rect 122 -70 123 -69
rect 123 -70 124 -69
rect 124 -70 125 -69
rect 125 -70 126 -69
rect 126 -70 127 -69
rect 127 -70 128 -69
rect 128 -70 129 -69
rect 129 -70 130 -69
rect 130 -70 131 -69
rect 131 -70 132 -69
rect 132 -70 133 -69
rect 133 -70 134 -69
rect 134 -70 135 -69
rect 135 -70 136 -69
rect 136 -70 137 -69
rect 137 -70 138 -69
rect 138 -70 139 -69
rect 139 -70 140 -69
rect 149 -70 150 -69
rect 150 -70 151 -69
rect 151 -70 152 -69
rect 152 -70 153 -69
rect 153 -70 154 -69
rect 154 -70 155 -69
rect 155 -70 156 -69
rect 156 -70 157 -69
rect 157 -70 158 -69
rect 158 -70 159 -69
rect 159 -70 160 -69
rect 160 -70 161 -69
rect 161 -70 162 -69
rect 162 -70 163 -69
rect 163 -70 164 -69
rect 164 -70 165 -69
rect 165 -70 166 -69
rect 166 -70 167 -69
rect 167 -70 168 -69
rect 168 -70 169 -69
rect 169 -70 170 -69
rect 170 -70 171 -69
rect 171 -70 172 -69
rect 181 -70 182 -69
rect 182 -70 183 -69
rect 183 -70 184 -69
rect 184 -70 185 -69
rect 185 -70 186 -69
rect 186 -70 187 -69
rect 187 -70 188 -69
rect 188 -70 189 -69
rect 189 -70 190 -69
rect 190 -70 191 -69
rect 191 -70 192 -69
rect 2 -71 3 -70
rect 3 -71 4 -70
rect 4 -71 5 -70
rect 5 -71 6 -70
rect 6 -71 7 -70
rect 7 -71 8 -70
rect 8 -71 9 -70
rect 9 -71 10 -70
rect 10 -71 11 -70
rect 11 -71 12 -70
rect 21 -71 22 -70
rect 22 -71 23 -70
rect 23 -71 24 -70
rect 24 -71 25 -70
rect 25 -71 26 -70
rect 26 -71 27 -70
rect 27 -71 28 -70
rect 28 -71 29 -70
rect 29 -71 30 -70
rect 30 -71 31 -70
rect 31 -71 32 -70
rect 32 -71 33 -70
rect 33 -71 34 -70
rect 34 -71 35 -70
rect 35 -71 36 -70
rect 36 -71 37 -70
rect 37 -71 38 -70
rect 38 -71 39 -70
rect 39 -71 40 -70
rect 40 -71 41 -70
rect 41 -71 42 -70
rect 42 -71 43 -70
rect 43 -71 44 -70
rect 53 -71 54 -70
rect 54 -71 55 -70
rect 55 -71 56 -70
rect 56 -71 57 -70
rect 57 -71 58 -70
rect 58 -71 59 -70
rect 59 -71 60 -70
rect 60 -71 61 -70
rect 61 -71 62 -70
rect 62 -71 63 -70
rect 63 -71 64 -70
rect 64 -71 65 -70
rect 65 -71 66 -70
rect 66 -71 67 -70
rect 67 -71 68 -70
rect 68 -71 69 -70
rect 69 -71 70 -70
rect 70 -71 71 -70
rect 71 -71 72 -70
rect 72 -71 73 -70
rect 73 -71 74 -70
rect 74 -71 75 -70
rect 75 -71 76 -70
rect 85 -71 86 -70
rect 86 -71 87 -70
rect 87 -71 88 -70
rect 88 -71 89 -70
rect 89 -71 90 -70
rect 90 -71 91 -70
rect 91 -71 92 -70
rect 92 -71 93 -70
rect 93 -71 94 -70
rect 94 -71 95 -70
rect 95 -71 96 -70
rect 96 -71 97 -70
rect 97 -71 98 -70
rect 98 -71 99 -70
rect 99 -71 100 -70
rect 100 -71 101 -70
rect 101 -71 102 -70
rect 102 -71 103 -70
rect 103 -71 104 -70
rect 104 -71 105 -70
rect 105 -71 106 -70
rect 106 -71 107 -70
rect 107 -71 108 -70
rect 117 -71 118 -70
rect 118 -71 119 -70
rect 119 -71 120 -70
rect 120 -71 121 -70
rect 121 -71 122 -70
rect 122 -71 123 -70
rect 123 -71 124 -70
rect 124 -71 125 -70
rect 125 -71 126 -70
rect 126 -71 127 -70
rect 127 -71 128 -70
rect 128 -71 129 -70
rect 129 -71 130 -70
rect 130 -71 131 -70
rect 131 -71 132 -70
rect 132 -71 133 -70
rect 133 -71 134 -70
rect 134 -71 135 -70
rect 135 -71 136 -70
rect 136 -71 137 -70
rect 137 -71 138 -70
rect 138 -71 139 -70
rect 139 -71 140 -70
rect 149 -71 150 -70
rect 150 -71 151 -70
rect 151 -71 152 -70
rect 152 -71 153 -70
rect 153 -71 154 -70
rect 154 -71 155 -70
rect 155 -71 156 -70
rect 156 -71 157 -70
rect 157 -71 158 -70
rect 158 -71 159 -70
rect 159 -71 160 -70
rect 160 -71 161 -70
rect 161 -71 162 -70
rect 162 -71 163 -70
rect 163 -71 164 -70
rect 164 -71 165 -70
rect 165 -71 166 -70
rect 166 -71 167 -70
rect 167 -71 168 -70
rect 168 -71 169 -70
rect 169 -71 170 -70
rect 170 -71 171 -70
rect 171 -71 172 -70
rect 181 -71 182 -70
rect 182 -71 183 -70
rect 183 -71 184 -70
rect 184 -71 185 -70
rect 185 -71 186 -70
rect 186 -71 187 -70
rect 187 -71 188 -70
rect 188 -71 189 -70
rect 189 -71 190 -70
rect 190 -71 191 -70
rect 191 -71 192 -70
rect 2 -72 3 -71
rect 3 -72 4 -71
rect 4 -72 5 -71
rect 5 -72 6 -71
rect 6 -72 7 -71
rect 7 -72 8 -71
rect 8 -72 9 -71
rect 9 -72 10 -71
rect 10 -72 11 -71
rect 11 -72 12 -71
rect 21 -72 22 -71
rect 22 -72 23 -71
rect 23 -72 24 -71
rect 24 -72 25 -71
rect 25 -72 26 -71
rect 26 -72 27 -71
rect 27 -72 28 -71
rect 28 -72 29 -71
rect 29 -72 30 -71
rect 30 -72 31 -71
rect 31 -72 32 -71
rect 32 -72 33 -71
rect 33 -72 34 -71
rect 34 -72 35 -71
rect 35 -72 36 -71
rect 36 -72 37 -71
rect 37 -72 38 -71
rect 38 -72 39 -71
rect 39 -72 40 -71
rect 40 -72 41 -71
rect 41 -72 42 -71
rect 42 -72 43 -71
rect 43 -72 44 -71
rect 53 -72 54 -71
rect 54 -72 55 -71
rect 55 -72 56 -71
rect 56 -72 57 -71
rect 57 -72 58 -71
rect 58 -72 59 -71
rect 59 -72 60 -71
rect 60 -72 61 -71
rect 61 -72 62 -71
rect 62 -72 63 -71
rect 63 -72 64 -71
rect 64 -72 65 -71
rect 65 -72 66 -71
rect 66 -72 67 -71
rect 67 -72 68 -71
rect 68 -72 69 -71
rect 69 -72 70 -71
rect 70 -72 71 -71
rect 71 -72 72 -71
rect 72 -72 73 -71
rect 73 -72 74 -71
rect 74 -72 75 -71
rect 75 -72 76 -71
rect 85 -72 86 -71
rect 86 -72 87 -71
rect 87 -72 88 -71
rect 88 -72 89 -71
rect 89 -72 90 -71
rect 90 -72 91 -71
rect 91 -72 92 -71
rect 92 -72 93 -71
rect 93 -72 94 -71
rect 94 -72 95 -71
rect 95 -72 96 -71
rect 96 -72 97 -71
rect 97 -72 98 -71
rect 98 -72 99 -71
rect 99 -72 100 -71
rect 100 -72 101 -71
rect 101 -72 102 -71
rect 102 -72 103 -71
rect 103 -72 104 -71
rect 104 -72 105 -71
rect 105 -72 106 -71
rect 106 -72 107 -71
rect 107 -72 108 -71
rect 117 -72 118 -71
rect 118 -72 119 -71
rect 119 -72 120 -71
rect 120 -72 121 -71
rect 121 -72 122 -71
rect 122 -72 123 -71
rect 123 -72 124 -71
rect 124 -72 125 -71
rect 125 -72 126 -71
rect 126 -72 127 -71
rect 127 -72 128 -71
rect 128 -72 129 -71
rect 129 -72 130 -71
rect 130 -72 131 -71
rect 131 -72 132 -71
rect 132 -72 133 -71
rect 133 -72 134 -71
rect 134 -72 135 -71
rect 135 -72 136 -71
rect 136 -72 137 -71
rect 137 -72 138 -71
rect 138 -72 139 -71
rect 139 -72 140 -71
rect 149 -72 150 -71
rect 150 -72 151 -71
rect 151 -72 152 -71
rect 152 -72 153 -71
rect 153 -72 154 -71
rect 154 -72 155 -71
rect 155 -72 156 -71
rect 156 -72 157 -71
rect 157 -72 158 -71
rect 158 -72 159 -71
rect 159 -72 160 -71
rect 160 -72 161 -71
rect 161 -72 162 -71
rect 162 -72 163 -71
rect 163 -72 164 -71
rect 164 -72 165 -71
rect 165 -72 166 -71
rect 166 -72 167 -71
rect 167 -72 168 -71
rect 168 -72 169 -71
rect 169 -72 170 -71
rect 170 -72 171 -71
rect 171 -72 172 -71
rect 181 -72 182 -71
rect 182 -72 183 -71
rect 183 -72 184 -71
rect 184 -72 185 -71
rect 185 -72 186 -71
rect 186 -72 187 -71
rect 187 -72 188 -71
rect 188 -72 189 -71
rect 189 -72 190 -71
rect 190 -72 191 -71
rect 191 -72 192 -71
rect 2 -73 3 -72
rect 3 -73 4 -72
rect 4 -73 5 -72
rect 5 -73 6 -72
rect 6 -73 7 -72
rect 7 -73 8 -72
rect 8 -73 9 -72
rect 9 -73 10 -72
rect 10 -73 11 -72
rect 11 -73 12 -72
rect 15 -73 16 -72
rect 16 -73 17 -72
rect 17 -73 18 -72
rect 21 -73 22 -72
rect 22 -73 23 -72
rect 23 -73 24 -72
rect 24 -73 25 -72
rect 25 -73 26 -72
rect 26 -73 27 -72
rect 27 -73 28 -72
rect 28 -73 29 -72
rect 29 -73 30 -72
rect 30 -73 31 -72
rect 31 -73 32 -72
rect 32 -73 33 -72
rect 33 -73 34 -72
rect 34 -73 35 -72
rect 35 -73 36 -72
rect 36 -73 37 -72
rect 37 -73 38 -72
rect 38 -73 39 -72
rect 39 -73 40 -72
rect 40 -73 41 -72
rect 41 -73 42 -72
rect 42 -73 43 -72
rect 43 -73 44 -72
rect 47 -73 48 -72
rect 48 -73 49 -72
rect 49 -73 50 -72
rect 53 -73 54 -72
rect 54 -73 55 -72
rect 55 -73 56 -72
rect 56 -73 57 -72
rect 57 -73 58 -72
rect 58 -73 59 -72
rect 59 -73 60 -72
rect 60 -73 61 -72
rect 61 -73 62 -72
rect 62 -73 63 -72
rect 63 -73 64 -72
rect 64 -73 65 -72
rect 65 -73 66 -72
rect 66 -73 67 -72
rect 67 -73 68 -72
rect 68 -73 69 -72
rect 69 -73 70 -72
rect 70 -73 71 -72
rect 71 -73 72 -72
rect 72 -73 73 -72
rect 73 -73 74 -72
rect 74 -73 75 -72
rect 75 -73 76 -72
rect 79 -73 80 -72
rect 80 -73 81 -72
rect 81 -73 82 -72
rect 85 -73 86 -72
rect 86 -73 87 -72
rect 87 -73 88 -72
rect 88 -73 89 -72
rect 89 -73 90 -72
rect 90 -73 91 -72
rect 91 -73 92 -72
rect 92 -73 93 -72
rect 93 -73 94 -72
rect 94 -73 95 -72
rect 95 -73 96 -72
rect 96 -73 97 -72
rect 97 -73 98 -72
rect 98 -73 99 -72
rect 99 -73 100 -72
rect 100 -73 101 -72
rect 101 -73 102 -72
rect 102 -73 103 -72
rect 103 -73 104 -72
rect 104 -73 105 -72
rect 105 -73 106 -72
rect 106 -73 107 -72
rect 107 -73 108 -72
rect 111 -73 112 -72
rect 112 -73 113 -72
rect 113 -73 114 -72
rect 117 -73 118 -72
rect 118 -73 119 -72
rect 119 -73 120 -72
rect 120 -73 121 -72
rect 121 -73 122 -72
rect 122 -73 123 -72
rect 123 -73 124 -72
rect 124 -73 125 -72
rect 125 -73 126 -72
rect 126 -73 127 -72
rect 127 -73 128 -72
rect 128 -73 129 -72
rect 129 -73 130 -72
rect 130 -73 131 -72
rect 131 -73 132 -72
rect 132 -73 133 -72
rect 133 -73 134 -72
rect 134 -73 135 -72
rect 135 -73 136 -72
rect 136 -73 137 -72
rect 137 -73 138 -72
rect 138 -73 139 -72
rect 139 -73 140 -72
rect 143 -73 144 -72
rect 144 -73 145 -72
rect 145 -73 146 -72
rect 149 -73 150 -72
rect 150 -73 151 -72
rect 151 -73 152 -72
rect 152 -73 153 -72
rect 153 -73 154 -72
rect 154 -73 155 -72
rect 155 -73 156 -72
rect 156 -73 157 -72
rect 157 -73 158 -72
rect 158 -73 159 -72
rect 159 -73 160 -72
rect 160 -73 161 -72
rect 161 -73 162 -72
rect 162 -73 163 -72
rect 163 -73 164 -72
rect 164 -73 165 -72
rect 165 -73 166 -72
rect 166 -73 167 -72
rect 167 -73 168 -72
rect 168 -73 169 -72
rect 169 -73 170 -72
rect 170 -73 171 -72
rect 171 -73 172 -72
rect 175 -73 176 -72
rect 176 -73 177 -72
rect 177 -73 178 -72
rect 181 -73 182 -72
rect 182 -73 183 -72
rect 183 -73 184 -72
rect 184 -73 185 -72
rect 185 -73 186 -72
rect 186 -73 187 -72
rect 187 -73 188 -72
rect 188 -73 189 -72
rect 189 -73 190 -72
rect 190 -73 191 -72
rect 191 -73 192 -72
rect 2 -74 3 -73
rect 3 -74 4 -73
rect 4 -74 5 -73
rect 5 -74 6 -73
rect 6 -74 7 -73
rect 7 -74 8 -73
rect 8 -74 9 -73
rect 9 -74 10 -73
rect 10 -74 11 -73
rect 11 -74 12 -73
rect 12 -74 13 -73
rect 14 -74 15 -73
rect 15 -74 16 -73
rect 16 -74 17 -73
rect 17 -74 18 -73
rect 18 -74 19 -73
rect 19 -74 20 -73
rect 20 -74 21 -73
rect 21 -74 22 -73
rect 22 -74 23 -73
rect 23 -74 24 -73
rect 24 -74 25 -73
rect 25 -74 26 -73
rect 26 -74 27 -73
rect 27 -74 28 -73
rect 28 -74 29 -73
rect 29 -74 30 -73
rect 30 -74 31 -73
rect 34 -74 35 -73
rect 35 -74 36 -73
rect 36 -74 37 -73
rect 37 -74 38 -73
rect 38 -74 39 -73
rect 39 -74 40 -73
rect 40 -74 41 -73
rect 41 -74 42 -73
rect 42 -74 43 -73
rect 43 -74 44 -73
rect 44 -74 45 -73
rect 46 -74 47 -73
rect 47 -74 48 -73
rect 48 -74 49 -73
rect 49 -74 50 -73
rect 50 -74 51 -73
rect 51 -74 52 -73
rect 52 -74 53 -73
rect 53 -74 54 -73
rect 54 -74 55 -73
rect 55 -74 56 -73
rect 56 -74 57 -73
rect 57 -74 58 -73
rect 58 -74 59 -73
rect 59 -74 60 -73
rect 60 -74 61 -73
rect 61 -74 62 -73
rect 62 -74 63 -73
rect 66 -74 67 -73
rect 67 -74 68 -73
rect 68 -74 69 -73
rect 69 -74 70 -73
rect 70 -74 71 -73
rect 71 -74 72 -73
rect 72 -74 73 -73
rect 73 -74 74 -73
rect 74 -74 75 -73
rect 75 -74 76 -73
rect 76 -74 77 -73
rect 78 -74 79 -73
rect 79 -74 80 -73
rect 80 -74 81 -73
rect 81 -74 82 -73
rect 82 -74 83 -73
rect 83 -74 84 -73
rect 84 -74 85 -73
rect 85 -74 86 -73
rect 86 -74 87 -73
rect 87 -74 88 -73
rect 88 -74 89 -73
rect 89 -74 90 -73
rect 90 -74 91 -73
rect 91 -74 92 -73
rect 92 -74 93 -73
rect 93 -74 94 -73
rect 94 -74 95 -73
rect 98 -74 99 -73
rect 99 -74 100 -73
rect 100 -74 101 -73
rect 101 -74 102 -73
rect 102 -74 103 -73
rect 103 -74 104 -73
rect 104 -74 105 -73
rect 105 -74 106 -73
rect 106 -74 107 -73
rect 107 -74 108 -73
rect 108 -74 109 -73
rect 110 -74 111 -73
rect 111 -74 112 -73
rect 112 -74 113 -73
rect 113 -74 114 -73
rect 114 -74 115 -73
rect 115 -74 116 -73
rect 116 -74 117 -73
rect 117 -74 118 -73
rect 118 -74 119 -73
rect 119 -74 120 -73
rect 120 -74 121 -73
rect 121 -74 122 -73
rect 122 -74 123 -73
rect 123 -74 124 -73
rect 124 -74 125 -73
rect 125 -74 126 -73
rect 126 -74 127 -73
rect 130 -74 131 -73
rect 131 -74 132 -73
rect 132 -74 133 -73
rect 133 -74 134 -73
rect 134 -74 135 -73
rect 135 -74 136 -73
rect 136 -74 137 -73
rect 137 -74 138 -73
rect 138 -74 139 -73
rect 139 -74 140 -73
rect 140 -74 141 -73
rect 142 -74 143 -73
rect 143 -74 144 -73
rect 144 -74 145 -73
rect 145 -74 146 -73
rect 146 -74 147 -73
rect 147 -74 148 -73
rect 148 -74 149 -73
rect 149 -74 150 -73
rect 150 -74 151 -73
rect 151 -74 152 -73
rect 152 -74 153 -73
rect 153 -74 154 -73
rect 154 -74 155 -73
rect 155 -74 156 -73
rect 156 -74 157 -73
rect 157 -74 158 -73
rect 158 -74 159 -73
rect 162 -74 163 -73
rect 163 -74 164 -73
rect 164 -74 165 -73
rect 165 -74 166 -73
rect 166 -74 167 -73
rect 167 -74 168 -73
rect 168 -74 169 -73
rect 169 -74 170 -73
rect 170 -74 171 -73
rect 171 -74 172 -73
rect 172 -74 173 -73
rect 174 -74 175 -73
rect 175 -74 176 -73
rect 176 -74 177 -73
rect 177 -74 178 -73
rect 178 -74 179 -73
rect 179 -74 180 -73
rect 180 -74 181 -73
rect 181 -74 182 -73
rect 182 -74 183 -73
rect 183 -74 184 -73
rect 184 -74 185 -73
rect 185 -74 186 -73
rect 186 -74 187 -73
rect 187 -74 188 -73
rect 188 -74 189 -73
rect 189 -74 190 -73
rect 190 -74 191 -73
rect 191 -74 192 -73
rect 2 -75 3 -74
rect 3 -75 4 -74
rect 4 -75 5 -74
rect 5 -75 6 -74
rect 6 -75 7 -74
rect 7 -75 8 -74
rect 8 -75 9 -74
rect 9 -75 10 -74
rect 10 -75 11 -74
rect 11 -75 12 -74
rect 12 -75 13 -74
rect 13 -75 14 -74
rect 14 -75 15 -74
rect 15 -75 16 -74
rect 16 -75 17 -74
rect 17 -75 18 -74
rect 18 -75 19 -74
rect 19 -75 20 -74
rect 20 -75 21 -74
rect 21 -75 22 -74
rect 22 -75 23 -74
rect 23 -75 24 -74
rect 24 -75 25 -74
rect 25 -75 26 -74
rect 26 -75 27 -74
rect 27 -75 28 -74
rect 28 -75 29 -74
rect 29 -75 30 -74
rect 30 -75 31 -74
rect 34 -75 35 -74
rect 35 -75 36 -74
rect 36 -75 37 -74
rect 37 -75 38 -74
rect 38 -75 39 -74
rect 39 -75 40 -74
rect 40 -75 41 -74
rect 41 -75 42 -74
rect 42 -75 43 -74
rect 43 -75 44 -74
rect 44 -75 45 -74
rect 45 -75 46 -74
rect 46 -75 47 -74
rect 47 -75 48 -74
rect 48 -75 49 -74
rect 49 -75 50 -74
rect 50 -75 51 -74
rect 51 -75 52 -74
rect 52 -75 53 -74
rect 53 -75 54 -74
rect 54 -75 55 -74
rect 55 -75 56 -74
rect 56 -75 57 -74
rect 57 -75 58 -74
rect 58 -75 59 -74
rect 59 -75 60 -74
rect 60 -75 61 -74
rect 61 -75 62 -74
rect 62 -75 63 -74
rect 66 -75 67 -74
rect 67 -75 68 -74
rect 68 -75 69 -74
rect 69 -75 70 -74
rect 70 -75 71 -74
rect 71 -75 72 -74
rect 72 -75 73 -74
rect 73 -75 74 -74
rect 74 -75 75 -74
rect 75 -75 76 -74
rect 76 -75 77 -74
rect 77 -75 78 -74
rect 78 -75 79 -74
rect 79 -75 80 -74
rect 80 -75 81 -74
rect 81 -75 82 -74
rect 82 -75 83 -74
rect 83 -75 84 -74
rect 84 -75 85 -74
rect 85 -75 86 -74
rect 86 -75 87 -74
rect 87 -75 88 -74
rect 88 -75 89 -74
rect 89 -75 90 -74
rect 90 -75 91 -74
rect 91 -75 92 -74
rect 92 -75 93 -74
rect 93 -75 94 -74
rect 94 -75 95 -74
rect 98 -75 99 -74
rect 99 -75 100 -74
rect 100 -75 101 -74
rect 101 -75 102 -74
rect 102 -75 103 -74
rect 103 -75 104 -74
rect 104 -75 105 -74
rect 105 -75 106 -74
rect 106 -75 107 -74
rect 107 -75 108 -74
rect 108 -75 109 -74
rect 109 -75 110 -74
rect 110 -75 111 -74
rect 111 -75 112 -74
rect 112 -75 113 -74
rect 113 -75 114 -74
rect 114 -75 115 -74
rect 115 -75 116 -74
rect 116 -75 117 -74
rect 117 -75 118 -74
rect 118 -75 119 -74
rect 119 -75 120 -74
rect 120 -75 121 -74
rect 121 -75 122 -74
rect 122 -75 123 -74
rect 123 -75 124 -74
rect 124 -75 125 -74
rect 125 -75 126 -74
rect 126 -75 127 -74
rect 130 -75 131 -74
rect 131 -75 132 -74
rect 132 -75 133 -74
rect 133 -75 134 -74
rect 134 -75 135 -74
rect 135 -75 136 -74
rect 136 -75 137 -74
rect 137 -75 138 -74
rect 138 -75 139 -74
rect 139 -75 140 -74
rect 140 -75 141 -74
rect 141 -75 142 -74
rect 142 -75 143 -74
rect 143 -75 144 -74
rect 144 -75 145 -74
rect 145 -75 146 -74
rect 146 -75 147 -74
rect 147 -75 148 -74
rect 148 -75 149 -74
rect 149 -75 150 -74
rect 150 -75 151 -74
rect 151 -75 152 -74
rect 152 -75 153 -74
rect 153 -75 154 -74
rect 154 -75 155 -74
rect 155 -75 156 -74
rect 156 -75 157 -74
rect 157 -75 158 -74
rect 158 -75 159 -74
rect 162 -75 163 -74
rect 163 -75 164 -74
rect 164 -75 165 -74
rect 165 -75 166 -74
rect 166 -75 167 -74
rect 167 -75 168 -74
rect 168 -75 169 -74
rect 169 -75 170 -74
rect 170 -75 171 -74
rect 171 -75 172 -74
rect 172 -75 173 -74
rect 173 -75 174 -74
rect 174 -75 175 -74
rect 175 -75 176 -74
rect 176 -75 177 -74
rect 177 -75 178 -74
rect 178 -75 179 -74
rect 179 -75 180 -74
rect 180 -75 181 -74
rect 181 -75 182 -74
rect 182 -75 183 -74
rect 183 -75 184 -74
rect 184 -75 185 -74
rect 185 -75 186 -74
rect 186 -75 187 -74
rect 187 -75 188 -74
rect 188 -75 189 -74
rect 189 -75 190 -74
rect 190 -75 191 -74
rect 191 -75 192 -74
rect 2 -76 3 -75
rect 3 -76 4 -75
rect 4 -76 5 -75
rect 5 -76 6 -75
rect 6 -76 7 -75
rect 7 -76 8 -75
rect 8 -76 9 -75
rect 9 -76 10 -75
rect 10 -76 11 -75
rect 11 -76 12 -75
rect 12 -76 13 -75
rect 13 -76 14 -75
rect 14 -76 15 -75
rect 15 -76 16 -75
rect 16 -76 17 -75
rect 17 -76 18 -75
rect 18 -76 19 -75
rect 19 -76 20 -75
rect 20 -76 21 -75
rect 21 -76 22 -75
rect 22 -76 23 -75
rect 23 -76 24 -75
rect 24 -76 25 -75
rect 25 -76 26 -75
rect 26 -76 27 -75
rect 27 -76 28 -75
rect 28 -76 29 -75
rect 29 -76 30 -75
rect 30 -76 31 -75
rect 35 -76 36 -75
rect 36 -76 37 -75
rect 37 -76 38 -75
rect 38 -76 39 -75
rect 39 -76 40 -75
rect 40 -76 41 -75
rect 41 -76 42 -75
rect 42 -76 43 -75
rect 43 -76 44 -75
rect 44 -76 45 -75
rect 45 -76 46 -75
rect 46 -76 47 -75
rect 47 -76 48 -75
rect 48 -76 49 -75
rect 49 -76 50 -75
rect 50 -76 51 -75
rect 51 -76 52 -75
rect 52 -76 53 -75
rect 53 -76 54 -75
rect 54 -76 55 -75
rect 55 -76 56 -75
rect 56 -76 57 -75
rect 57 -76 58 -75
rect 58 -76 59 -75
rect 59 -76 60 -75
rect 60 -76 61 -75
rect 61 -76 62 -75
rect 62 -76 63 -75
rect 67 -76 68 -75
rect 68 -76 69 -75
rect 69 -76 70 -75
rect 70 -76 71 -75
rect 71 -76 72 -75
rect 72 -76 73 -75
rect 73 -76 74 -75
rect 74 -76 75 -75
rect 75 -76 76 -75
rect 76 -76 77 -75
rect 77 -76 78 -75
rect 78 -76 79 -75
rect 79 -76 80 -75
rect 80 -76 81 -75
rect 81 -76 82 -75
rect 82 -76 83 -75
rect 83 -76 84 -75
rect 84 -76 85 -75
rect 85 -76 86 -75
rect 86 -76 87 -75
rect 87 -76 88 -75
rect 88 -76 89 -75
rect 89 -76 90 -75
rect 90 -76 91 -75
rect 91 -76 92 -75
rect 92 -76 93 -75
rect 93 -76 94 -75
rect 94 -76 95 -75
rect 99 -76 100 -75
rect 100 -76 101 -75
rect 101 -76 102 -75
rect 102 -76 103 -75
rect 103 -76 104 -75
rect 104 -76 105 -75
rect 105 -76 106 -75
rect 106 -76 107 -75
rect 107 -76 108 -75
rect 108 -76 109 -75
rect 109 -76 110 -75
rect 110 -76 111 -75
rect 111 -76 112 -75
rect 112 -76 113 -75
rect 113 -76 114 -75
rect 114 -76 115 -75
rect 115 -76 116 -75
rect 116 -76 117 -75
rect 117 -76 118 -75
rect 118 -76 119 -75
rect 119 -76 120 -75
rect 120 -76 121 -75
rect 121 -76 122 -75
rect 122 -76 123 -75
rect 123 -76 124 -75
rect 124 -76 125 -75
rect 125 -76 126 -75
rect 126 -76 127 -75
rect 131 -76 132 -75
rect 132 -76 133 -75
rect 133 -76 134 -75
rect 134 -76 135 -75
rect 135 -76 136 -75
rect 136 -76 137 -75
rect 137 -76 138 -75
rect 138 -76 139 -75
rect 139 -76 140 -75
rect 140 -76 141 -75
rect 141 -76 142 -75
rect 142 -76 143 -75
rect 143 -76 144 -75
rect 144 -76 145 -75
rect 145 -76 146 -75
rect 146 -76 147 -75
rect 147 -76 148 -75
rect 148 -76 149 -75
rect 149 -76 150 -75
rect 150 -76 151 -75
rect 151 -76 152 -75
rect 152 -76 153 -75
rect 153 -76 154 -75
rect 154 -76 155 -75
rect 155 -76 156 -75
rect 156 -76 157 -75
rect 157 -76 158 -75
rect 158 -76 159 -75
rect 163 -76 164 -75
rect 164 -76 165 -75
rect 165 -76 166 -75
rect 166 -76 167 -75
rect 167 -76 168 -75
rect 168 -76 169 -75
rect 169 -76 170 -75
rect 170 -76 171 -75
rect 171 -76 172 -75
rect 172 -76 173 -75
rect 173 -76 174 -75
rect 174 -76 175 -75
rect 175 -76 176 -75
rect 176 -76 177 -75
rect 177 -76 178 -75
rect 178 -76 179 -75
rect 179 -76 180 -75
rect 180 -76 181 -75
rect 181 -76 182 -75
rect 182 -76 183 -75
rect 183 -76 184 -75
rect 184 -76 185 -75
rect 185 -76 186 -75
rect 186 -76 187 -75
rect 187 -76 188 -75
rect 188 -76 189 -75
rect 189 -76 190 -75
rect 190 -76 191 -75
rect 191 -76 192 -75
rect 2 -77 3 -76
rect 3 -77 4 -76
rect 4 -77 5 -76
rect 5 -77 6 -76
rect 6 -77 7 -76
rect 7 -77 8 -76
rect 8 -77 9 -76
rect 9 -77 10 -76
rect 10 -77 11 -76
rect 11 -77 12 -76
rect 12 -77 13 -76
rect 13 -77 14 -76
rect 14 -77 15 -76
rect 15 -77 16 -76
rect 16 -77 17 -76
rect 17 -77 18 -76
rect 18 -77 19 -76
rect 19 -77 20 -76
rect 20 -77 21 -76
rect 21 -77 22 -76
rect 22 -77 23 -76
rect 23 -77 24 -76
rect 24 -77 25 -76
rect 25 -77 26 -76
rect 26 -77 27 -76
rect 27 -77 28 -76
rect 28 -77 29 -76
rect 29 -77 30 -76
rect 30 -77 31 -76
rect 35 -77 36 -76
rect 36 -77 37 -76
rect 37 -77 38 -76
rect 38 -77 39 -76
rect 39 -77 40 -76
rect 40 -77 41 -76
rect 41 -77 42 -76
rect 42 -77 43 -76
rect 43 -77 44 -76
rect 44 -77 45 -76
rect 45 -77 46 -76
rect 46 -77 47 -76
rect 47 -77 48 -76
rect 48 -77 49 -76
rect 49 -77 50 -76
rect 50 -77 51 -76
rect 51 -77 52 -76
rect 52 -77 53 -76
rect 53 -77 54 -76
rect 54 -77 55 -76
rect 55 -77 56 -76
rect 56 -77 57 -76
rect 57 -77 58 -76
rect 58 -77 59 -76
rect 59 -77 60 -76
rect 60 -77 61 -76
rect 61 -77 62 -76
rect 67 -77 68 -76
rect 68 -77 69 -76
rect 69 -77 70 -76
rect 70 -77 71 -76
rect 71 -77 72 -76
rect 72 -77 73 -76
rect 73 -77 74 -76
rect 74 -77 75 -76
rect 75 -77 76 -76
rect 76 -77 77 -76
rect 77 -77 78 -76
rect 78 -77 79 -76
rect 79 -77 80 -76
rect 80 -77 81 -76
rect 81 -77 82 -76
rect 82 -77 83 -76
rect 83 -77 84 -76
rect 84 -77 85 -76
rect 85 -77 86 -76
rect 86 -77 87 -76
rect 87 -77 88 -76
rect 88 -77 89 -76
rect 89 -77 90 -76
rect 90 -77 91 -76
rect 91 -77 92 -76
rect 92 -77 93 -76
rect 93 -77 94 -76
rect 94 -77 95 -76
rect 99 -77 100 -76
rect 100 -77 101 -76
rect 101 -77 102 -76
rect 102 -77 103 -76
rect 103 -77 104 -76
rect 104 -77 105 -76
rect 105 -77 106 -76
rect 106 -77 107 -76
rect 107 -77 108 -76
rect 108 -77 109 -76
rect 109 -77 110 -76
rect 110 -77 111 -76
rect 111 -77 112 -76
rect 112 -77 113 -76
rect 113 -77 114 -76
rect 114 -77 115 -76
rect 115 -77 116 -76
rect 116 -77 117 -76
rect 117 -77 118 -76
rect 118 -77 119 -76
rect 119 -77 120 -76
rect 120 -77 121 -76
rect 121 -77 122 -76
rect 122 -77 123 -76
rect 123 -77 124 -76
rect 124 -77 125 -76
rect 125 -77 126 -76
rect 131 -77 132 -76
rect 132 -77 133 -76
rect 133 -77 134 -76
rect 134 -77 135 -76
rect 135 -77 136 -76
rect 136 -77 137 -76
rect 137 -77 138 -76
rect 138 -77 139 -76
rect 139 -77 140 -76
rect 140 -77 141 -76
rect 141 -77 142 -76
rect 142 -77 143 -76
rect 143 -77 144 -76
rect 144 -77 145 -76
rect 145 -77 146 -76
rect 146 -77 147 -76
rect 147 -77 148 -76
rect 148 -77 149 -76
rect 149 -77 150 -76
rect 150 -77 151 -76
rect 151 -77 152 -76
rect 152 -77 153 -76
rect 153 -77 154 -76
rect 154 -77 155 -76
rect 155 -77 156 -76
rect 156 -77 157 -76
rect 157 -77 158 -76
rect 158 -77 159 -76
rect 163 -77 164 -76
rect 164 -77 165 -76
rect 165 -77 166 -76
rect 166 -77 167 -76
rect 167 -77 168 -76
rect 168 -77 169 -76
rect 169 -77 170 -76
rect 170 -77 171 -76
rect 171 -77 172 -76
rect 172 -77 173 -76
rect 173 -77 174 -76
rect 174 -77 175 -76
rect 175 -77 176 -76
rect 176 -77 177 -76
rect 177 -77 178 -76
rect 178 -77 179 -76
rect 179 -77 180 -76
rect 180 -77 181 -76
rect 181 -77 182 -76
rect 182 -77 183 -76
rect 183 -77 184 -76
rect 184 -77 185 -76
rect 185 -77 186 -76
rect 186 -77 187 -76
rect 187 -77 188 -76
rect 188 -77 189 -76
rect 189 -77 190 -76
rect 190 -77 191 -76
rect 191 -77 192 -76
rect 2 -78 3 -77
rect 3 -78 4 -77
rect 4 -78 5 -77
rect 5 -78 6 -77
rect 6 -78 7 -77
rect 7 -78 8 -77
rect 8 -78 9 -77
rect 9 -78 10 -77
rect 10 -78 11 -77
rect 11 -78 12 -77
rect 12 -78 13 -77
rect 13 -78 14 -77
rect 14 -78 15 -77
rect 15 -78 16 -77
rect 16 -78 17 -77
rect 17 -78 18 -77
rect 18 -78 19 -77
rect 19 -78 20 -77
rect 20 -78 21 -77
rect 21 -78 22 -77
rect 22 -78 23 -77
rect 23 -78 24 -77
rect 24 -78 25 -77
rect 26 -78 27 -77
rect 27 -78 28 -77
rect 28 -78 29 -77
rect 37 -78 38 -77
rect 38 -78 39 -77
rect 41 -78 42 -77
rect 42 -78 43 -77
rect 43 -78 44 -77
rect 44 -78 45 -77
rect 45 -78 46 -77
rect 46 -78 47 -77
rect 47 -78 48 -77
rect 48 -78 49 -77
rect 49 -78 50 -77
rect 50 -78 51 -77
rect 51 -78 52 -77
rect 52 -78 53 -77
rect 53 -78 54 -77
rect 54 -78 55 -77
rect 55 -78 56 -77
rect 56 -78 57 -77
rect 58 -78 59 -77
rect 59 -78 60 -77
rect 60 -78 61 -77
rect 68 -78 69 -77
rect 69 -78 70 -77
rect 70 -78 71 -77
rect 73 -78 74 -77
rect 74 -78 75 -77
rect 75 -78 76 -77
rect 76 -78 77 -77
rect 77 -78 78 -77
rect 78 -78 79 -77
rect 79 -78 80 -77
rect 80 -78 81 -77
rect 81 -78 82 -77
rect 82 -78 83 -77
rect 83 -78 84 -77
rect 84 -78 85 -77
rect 85 -78 86 -77
rect 86 -78 87 -77
rect 87 -78 88 -77
rect 88 -78 89 -77
rect 90 -78 91 -77
rect 91 -78 92 -77
rect 92 -78 93 -77
rect 101 -78 102 -77
rect 102 -78 103 -77
rect 105 -78 106 -77
rect 106 -78 107 -77
rect 107 -78 108 -77
rect 108 -78 109 -77
rect 109 -78 110 -77
rect 110 -78 111 -77
rect 111 -78 112 -77
rect 112 -78 113 -77
rect 113 -78 114 -77
rect 114 -78 115 -77
rect 115 -78 116 -77
rect 116 -78 117 -77
rect 117 -78 118 -77
rect 118 -78 119 -77
rect 119 -78 120 -77
rect 120 -78 121 -77
rect 122 -78 123 -77
rect 123 -78 124 -77
rect 124 -78 125 -77
rect 132 -78 133 -77
rect 133 -78 134 -77
rect 134 -78 135 -77
rect 137 -78 138 -77
rect 138 -78 139 -77
rect 139 -78 140 -77
rect 140 -78 141 -77
rect 141 -78 142 -77
rect 142 -78 143 -77
rect 143 -78 144 -77
rect 144 -78 145 -77
rect 145 -78 146 -77
rect 146 -78 147 -77
rect 147 -78 148 -77
rect 148 -78 149 -77
rect 149 -78 150 -77
rect 150 -78 151 -77
rect 151 -78 152 -77
rect 152 -78 153 -77
rect 154 -78 155 -77
rect 155 -78 156 -77
rect 156 -78 157 -77
rect 165 -78 166 -77
rect 166 -78 167 -77
rect 169 -78 170 -77
rect 170 -78 171 -77
rect 171 -78 172 -77
rect 172 -78 173 -77
rect 173 -78 174 -77
rect 174 -78 175 -77
rect 175 -78 176 -77
rect 176 -78 177 -77
rect 177 -78 178 -77
rect 178 -78 179 -77
rect 179 -78 180 -77
rect 180 -78 181 -77
rect 181 -78 182 -77
rect 182 -78 183 -77
rect 183 -78 184 -77
rect 184 -78 185 -77
rect 185 -78 186 -77
rect 186 -78 187 -77
rect 187 -78 188 -77
rect 188 -78 189 -77
rect 189 -78 190 -77
rect 190 -78 191 -77
rect 191 -78 192 -77
rect 2 -79 3 -78
rect 3 -79 4 -78
rect 4 -79 5 -78
rect 5 -79 6 -78
rect 6 -79 7 -78
rect 7 -79 8 -78
rect 8 -79 9 -78
rect 9 -79 10 -78
rect 10 -79 11 -78
rect 11 -79 12 -78
rect 12 -79 13 -78
rect 13 -79 14 -78
rect 14 -79 15 -78
rect 15 -79 16 -78
rect 16 -79 17 -78
rect 17 -79 18 -78
rect 18 -79 19 -78
rect 19 -79 20 -78
rect 20 -79 21 -78
rect 21 -79 22 -78
rect 22 -79 23 -78
rect 23 -79 24 -78
rect 24 -79 25 -78
rect 41 -79 42 -78
rect 42 -79 43 -78
rect 43 -79 44 -78
rect 44 -79 45 -78
rect 45 -79 46 -78
rect 46 -79 47 -78
rect 47 -79 48 -78
rect 48 -79 49 -78
rect 49 -79 50 -78
rect 50 -79 51 -78
rect 51 -79 52 -78
rect 52 -79 53 -78
rect 53 -79 54 -78
rect 54 -79 55 -78
rect 55 -79 56 -78
rect 56 -79 57 -78
rect 73 -79 74 -78
rect 74 -79 75 -78
rect 75 -79 76 -78
rect 76 -79 77 -78
rect 77 -79 78 -78
rect 78 -79 79 -78
rect 79 -79 80 -78
rect 80 -79 81 -78
rect 81 -79 82 -78
rect 82 -79 83 -78
rect 83 -79 84 -78
rect 84 -79 85 -78
rect 85 -79 86 -78
rect 86 -79 87 -78
rect 87 -79 88 -78
rect 88 -79 89 -78
rect 105 -79 106 -78
rect 106 -79 107 -78
rect 107 -79 108 -78
rect 108 -79 109 -78
rect 109 -79 110 -78
rect 110 -79 111 -78
rect 111 -79 112 -78
rect 112 -79 113 -78
rect 113 -79 114 -78
rect 114 -79 115 -78
rect 115 -79 116 -78
rect 116 -79 117 -78
rect 117 -79 118 -78
rect 118 -79 119 -78
rect 119 -79 120 -78
rect 120 -79 121 -78
rect 137 -79 138 -78
rect 138 -79 139 -78
rect 139 -79 140 -78
rect 140 -79 141 -78
rect 141 -79 142 -78
rect 142 -79 143 -78
rect 143 -79 144 -78
rect 144 -79 145 -78
rect 145 -79 146 -78
rect 146 -79 147 -78
rect 147 -79 148 -78
rect 148 -79 149 -78
rect 149 -79 150 -78
rect 150 -79 151 -78
rect 151 -79 152 -78
rect 152 -79 153 -78
rect 169 -79 170 -78
rect 170 -79 171 -78
rect 171 -79 172 -78
rect 172 -79 173 -78
rect 173 -79 174 -78
rect 174 -79 175 -78
rect 175 -79 176 -78
rect 176 -79 177 -78
rect 177 -79 178 -78
rect 178 -79 179 -78
rect 179 -79 180 -78
rect 180 -79 181 -78
rect 181 -79 182 -78
rect 182 -79 183 -78
rect 183 -79 184 -78
rect 184 -79 185 -78
rect 185 -79 186 -78
rect 186 -79 187 -78
rect 187 -79 188 -78
rect 188 -79 189 -78
rect 189 -79 190 -78
rect 190 -79 191 -78
rect 191 -79 192 -78
rect 192 -79 193 -78
rect 193 -79 194 -78
rect 194 -79 195 -78
rect 195 -79 196 -78
rect 196 -79 197 -78
rect 197 -79 198 -78
rect 198 -79 199 -78
rect 199 -79 200 -78
rect 200 -79 201 -78
rect 201 -79 202 -78
rect 202 -79 203 -78
rect 203 -79 204 -78
rect 204 -79 205 -78
rect 205 -79 206 -78
rect 206 -79 207 -78
rect 207 -79 208 -78
rect 208 -79 209 -78
rect 209 -79 210 -78
rect 210 -79 211 -78
rect 211 -79 212 -78
rect 212 -79 213 -78
rect 213 -79 214 -78
rect 214 -79 215 -78
rect 215 -79 216 -78
rect 216 -79 217 -78
rect 217 -79 218 -78
rect 218 -79 219 -78
rect 219 -79 220 -78
rect 220 -79 221 -78
rect 221 -79 222 -78
rect 222 -79 223 -78
rect 223 -79 224 -78
rect 224 -79 225 -78
rect 225 -79 226 -78
rect 226 -79 227 -78
rect 227 -79 228 -78
rect 228 -79 229 -78
rect 229 -79 230 -78
rect 230 -79 231 -78
rect 231 -79 232 -78
rect 232 -79 233 -78
rect 233 -79 234 -78
rect 234 -79 235 -78
rect 235 -79 236 -78
rect 236 -79 237 -78
rect 237 -79 238 -78
rect 238 -79 239 -78
rect 239 -79 240 -78
rect 240 -79 241 -78
rect 241 -79 242 -78
rect 242 -79 243 -78
rect 243 -79 244 -78
rect 244 -79 245 -78
rect 245 -79 246 -78
rect 246 -79 247 -78
rect 247 -79 248 -78
rect 248 -79 249 -78
rect 249 -79 250 -78
rect 250 -79 251 -78
rect 251 -79 252 -78
rect 252 -79 253 -78
rect 253 -79 254 -78
rect 254 -79 255 -78
rect 255 -79 256 -78
rect 256 -79 257 -78
rect 257 -79 258 -78
rect 258 -79 259 -78
rect 259 -79 260 -78
rect 260 -79 261 -78
rect 261 -79 262 -78
rect 262 -79 263 -78
rect 263 -79 264 -78
rect 264 -79 265 -78
rect 265 -79 266 -78
rect 266 -79 267 -78
rect 267 -79 268 -78
rect 268 -79 269 -78
rect 269 -79 270 -78
rect 270 -79 271 -78
rect 271 -79 272 -78
rect 272 -79 273 -78
rect 273 -79 274 -78
rect 274 -79 275 -78
rect 275 -79 276 -78
rect 276 -79 277 -78
rect 277 -79 278 -78
rect 278 -79 279 -78
rect 279 -79 280 -78
rect 280 -79 281 -78
rect 281 -79 282 -78
rect 282 -79 283 -78
rect 283 -79 284 -78
rect 284 -79 285 -78
rect 285 -79 286 -78
rect 286 -79 287 -78
rect 287 -79 288 -78
rect 288 -79 289 -78
rect 289 -79 290 -78
rect 290 -79 291 -78
rect 291 -79 292 -78
rect 292 -79 293 -78
rect 293 -79 294 -78
rect 294 -79 295 -78
rect 295 -79 296 -78
rect 296 -79 297 -78
rect 297 -79 298 -78
rect 298 -79 299 -78
rect 299 -79 300 -78
rect 300 -79 301 -78
rect 301 -79 302 -78
rect 302 -79 303 -78
rect 303 -79 304 -78
rect 304 -79 305 -78
rect 305 -79 306 -78
rect 306 -79 307 -78
rect 307 -79 308 -78
rect 308 -79 309 -78
rect 309 -79 310 -78
rect 310 -79 311 -78
rect 311 -79 312 -78
rect 312 -79 313 -78
rect 313 -79 314 -78
rect 314 -79 315 -78
rect 315 -79 316 -78
rect 316 -79 317 -78
rect 317 -79 318 -78
rect 318 -79 319 -78
rect 319 -79 320 -78
rect 320 -79 321 -78
rect 321 -79 322 -78
rect 322 -79 323 -78
rect 323 -79 324 -78
rect 324 -79 325 -78
rect 325 -79 326 -78
rect 326 -79 327 -78
rect 327 -79 328 -78
rect 328 -79 329 -78
rect 329 -79 330 -78
rect 330 -79 331 -78
rect 331 -79 332 -78
rect 332 -79 333 -78
rect 333 -79 334 -78
rect 334 -79 335 -78
rect 335 -79 336 -78
rect 336 -79 337 -78
rect 337 -79 338 -78
rect 338 -79 339 -78
rect 339 -79 340 -78
rect 340 -79 341 -78
rect 341 -79 342 -78
rect 342 -79 343 -78
rect 343 -79 344 -78
rect 344 -79 345 -78
rect 345 -79 346 -78
rect 346 -79 347 -78
rect 347 -79 348 -78
rect 348 -79 349 -78
rect 349 -79 350 -78
rect 350 -79 351 -78
rect 351 -79 352 -78
rect 352 -79 353 -78
rect 353 -79 354 -78
rect 354 -79 355 -78
rect 355 -79 356 -78
rect 356 -79 357 -78
rect 357 -79 358 -78
rect 358 -79 359 -78
rect 359 -79 360 -78
rect 360 -79 361 -78
rect 361 -79 362 -78
rect 362 -79 363 -78
rect 363 -79 364 -78
rect 364 -79 365 -78
rect 365 -79 366 -78
rect 366 -79 367 -78
rect 367 -79 368 -78
rect 368 -79 369 -78
rect 369 -79 370 -78
rect 370 -79 371 -78
rect 371 -79 372 -78
rect 372 -79 373 -78
rect 373 -79 374 -78
rect 374 -79 375 -78
rect 375 -79 376 -78
rect 376 -79 377 -78
rect 377 -79 378 -78
rect 378 -79 379 -78
rect 379 -79 380 -78
rect 380 -79 381 -78
rect 381 -79 382 -78
rect 382 -79 383 -78
rect 383 -79 384 -78
rect 384 -79 385 -78
rect 385 -79 386 -78
rect 386 -79 387 -78
rect 387 -79 388 -78
rect 388 -79 389 -78
rect 389 -79 390 -78
rect 390 -79 391 -78
rect 391 -79 392 -78
rect 392 -79 393 -78
rect 393 -79 394 -78
rect 394 -79 395 -78
rect 395 -79 396 -78
rect 396 -79 397 -78
rect 397 -79 398 -78
rect 398 -79 399 -78
rect 399 -79 400 -78
rect 400 -79 401 -78
rect 401 -79 402 -78
rect 402 -79 403 -78
rect 403 -79 404 -78
rect 404 -79 405 -78
rect 405 -79 406 -78
rect 406 -79 407 -78
rect 407 -79 408 -78
rect 408 -79 409 -78
rect 409 -79 410 -78
rect 410 -79 411 -78
rect 411 -79 412 -78
rect 412 -79 413 -78
rect 413 -79 414 -78
rect 414 -79 415 -78
rect 415 -79 416 -78
rect 416 -79 417 -78
rect 417 -79 418 -78
rect 418 -79 419 -78
rect 419 -79 420 -78
rect 420 -79 421 -78
rect 421 -79 422 -78
rect 422 -79 423 -78
rect 423 -79 424 -78
rect 424 -79 425 -78
rect 425 -79 426 -78
rect 426 -79 427 -78
rect 427 -79 428 -78
rect 428 -79 429 -78
rect 429 -79 430 -78
rect 430 -79 431 -78
rect 431 -79 432 -78
rect 432 -79 433 -78
rect 433 -79 434 -78
rect 434 -79 435 -78
rect 435 -79 436 -78
rect 436 -79 437 -78
rect 437 -79 438 -78
rect 438 -79 439 -78
rect 439 -79 440 -78
rect 440 -79 441 -78
rect 441 -79 442 -78
rect 442 -79 443 -78
rect 443 -79 444 -78
rect 444 -79 445 -78
rect 445 -79 446 -78
rect 446 -79 447 -78
rect 447 -79 448 -78
rect 448 -79 449 -78
rect 449 -79 450 -78
rect 450 -79 451 -78
rect 451 -79 452 -78
rect 452 -79 453 -78
rect 453 -79 454 -78
rect 454 -79 455 -78
rect 455 -79 456 -78
rect 456 -79 457 -78
rect 457 -79 458 -78
rect 458 -79 459 -78
rect 459 -79 460 -78
rect 460 -79 461 -78
rect 461 -79 462 -78
rect 462 -79 463 -78
rect 463 -79 464 -78
rect 464 -79 465 -78
rect 465 -79 466 -78
rect 466 -79 467 -78
rect 467 -79 468 -78
rect 468 -79 469 -78
rect 469 -79 470 -78
rect 470 -79 471 -78
rect 471 -79 472 -78
rect 472 -79 473 -78
rect 473 -79 474 -78
rect 474 -79 475 -78
rect 475 -79 476 -78
rect 476 -79 477 -78
rect 477 -79 478 -78
rect 478 -79 479 -78
rect 479 -79 480 -78
rect 2 -80 3 -79
rect 3 -80 4 -79
rect 4 -80 5 -79
rect 5 -80 6 -79
rect 6 -80 7 -79
rect 7 -80 8 -79
rect 8 -80 9 -79
rect 9 -80 10 -79
rect 10 -80 11 -79
rect 11 -80 12 -79
rect 12 -80 13 -79
rect 13 -80 14 -79
rect 14 -80 15 -79
rect 15 -80 16 -79
rect 16 -80 17 -79
rect 17 -80 18 -79
rect 18 -80 19 -79
rect 19 -80 20 -79
rect 20 -80 21 -79
rect 21 -80 22 -79
rect 22 -80 23 -79
rect 23 -80 24 -79
rect 24 -80 25 -79
rect 41 -80 42 -79
rect 42 -80 43 -79
rect 43 -80 44 -79
rect 44 -80 45 -79
rect 45 -80 46 -79
rect 46 -80 47 -79
rect 47 -80 48 -79
rect 48 -80 49 -79
rect 49 -80 50 -79
rect 50 -80 51 -79
rect 51 -80 52 -79
rect 52 -80 53 -79
rect 53 -80 54 -79
rect 54 -80 55 -79
rect 55 -80 56 -79
rect 56 -80 57 -79
rect 73 -80 74 -79
rect 74 -80 75 -79
rect 75 -80 76 -79
rect 76 -80 77 -79
rect 77 -80 78 -79
rect 78 -80 79 -79
rect 79 -80 80 -79
rect 80 -80 81 -79
rect 81 -80 82 -79
rect 82 -80 83 -79
rect 83 -80 84 -79
rect 84 -80 85 -79
rect 85 -80 86 -79
rect 86 -80 87 -79
rect 87 -80 88 -79
rect 88 -80 89 -79
rect 105 -80 106 -79
rect 106 -80 107 -79
rect 107 -80 108 -79
rect 108 -80 109 -79
rect 109 -80 110 -79
rect 110 -80 111 -79
rect 111 -80 112 -79
rect 112 -80 113 -79
rect 113 -80 114 -79
rect 114 -80 115 -79
rect 115 -80 116 -79
rect 116 -80 117 -79
rect 117 -80 118 -79
rect 118 -80 119 -79
rect 119 -80 120 -79
rect 120 -80 121 -79
rect 137 -80 138 -79
rect 138 -80 139 -79
rect 139 -80 140 -79
rect 140 -80 141 -79
rect 141 -80 142 -79
rect 142 -80 143 -79
rect 143 -80 144 -79
rect 144 -80 145 -79
rect 145 -80 146 -79
rect 146 -80 147 -79
rect 147 -80 148 -79
rect 148 -80 149 -79
rect 149 -80 150 -79
rect 150 -80 151 -79
rect 151 -80 152 -79
rect 152 -80 153 -79
rect 169 -80 170 -79
rect 170 -80 171 -79
rect 171 -80 172 -79
rect 172 -80 173 -79
rect 173 -80 174 -79
rect 174 -80 175 -79
rect 175 -80 176 -79
rect 176 -80 177 -79
rect 177 -80 178 -79
rect 178 -80 179 -79
rect 179 -80 180 -79
rect 180 -80 181 -79
rect 181 -80 182 -79
rect 182 -80 183 -79
rect 183 -80 184 -79
rect 184 -80 185 -79
rect 185 -80 186 -79
rect 186 -80 187 -79
rect 187 -80 188 -79
rect 188 -80 189 -79
rect 189 -80 190 -79
rect 190 -80 191 -79
rect 191 -80 192 -79
rect 192 -80 193 -79
rect 193 -80 194 -79
rect 194 -80 195 -79
rect 195 -80 196 -79
rect 196 -80 197 -79
rect 197 -80 198 -79
rect 198 -80 199 -79
rect 199 -80 200 -79
rect 200 -80 201 -79
rect 201 -80 202 -79
rect 202 -80 203 -79
rect 203 -80 204 -79
rect 204 -80 205 -79
rect 205 -80 206 -79
rect 206 -80 207 -79
rect 207 -80 208 -79
rect 208 -80 209 -79
rect 209 -80 210 -79
rect 210 -80 211 -79
rect 211 -80 212 -79
rect 212 -80 213 -79
rect 213 -80 214 -79
rect 214 -80 215 -79
rect 215 -80 216 -79
rect 216 -80 217 -79
rect 217 -80 218 -79
rect 218 -80 219 -79
rect 219 -80 220 -79
rect 220 -80 221 -79
rect 221 -80 222 -79
rect 222 -80 223 -79
rect 223 -80 224 -79
rect 224 -80 225 -79
rect 225 -80 226 -79
rect 226 -80 227 -79
rect 227 -80 228 -79
rect 228 -80 229 -79
rect 229 -80 230 -79
rect 230 -80 231 -79
rect 231 -80 232 -79
rect 232 -80 233 -79
rect 233 -80 234 -79
rect 234 -80 235 -79
rect 235 -80 236 -79
rect 236 -80 237 -79
rect 237 -80 238 -79
rect 238 -80 239 -79
rect 239 -80 240 -79
rect 240 -80 241 -79
rect 241 -80 242 -79
rect 242 -80 243 -79
rect 243 -80 244 -79
rect 244 -80 245 -79
rect 245 -80 246 -79
rect 246 -80 247 -79
rect 247 -80 248 -79
rect 248 -80 249 -79
rect 249 -80 250 -79
rect 250 -80 251 -79
rect 251 -80 252 -79
rect 252 -80 253 -79
rect 253 -80 254 -79
rect 254 -80 255 -79
rect 255 -80 256 -79
rect 256 -80 257 -79
rect 257 -80 258 -79
rect 258 -80 259 -79
rect 259 -80 260 -79
rect 260 -80 261 -79
rect 261 -80 262 -79
rect 262 -80 263 -79
rect 263 -80 264 -79
rect 264 -80 265 -79
rect 265 -80 266 -79
rect 266 -80 267 -79
rect 267 -80 268 -79
rect 268 -80 269 -79
rect 269 -80 270 -79
rect 270 -80 271 -79
rect 271 -80 272 -79
rect 272 -80 273 -79
rect 273 -80 274 -79
rect 274 -80 275 -79
rect 275 -80 276 -79
rect 276 -80 277 -79
rect 277 -80 278 -79
rect 278 -80 279 -79
rect 279 -80 280 -79
rect 280 -80 281 -79
rect 281 -80 282 -79
rect 282 -80 283 -79
rect 283 -80 284 -79
rect 284 -80 285 -79
rect 285 -80 286 -79
rect 286 -80 287 -79
rect 287 -80 288 -79
rect 288 -80 289 -79
rect 289 -80 290 -79
rect 290 -80 291 -79
rect 291 -80 292 -79
rect 292 -80 293 -79
rect 293 -80 294 -79
rect 294 -80 295 -79
rect 295 -80 296 -79
rect 296 -80 297 -79
rect 297 -80 298 -79
rect 298 -80 299 -79
rect 299 -80 300 -79
rect 300 -80 301 -79
rect 301 -80 302 -79
rect 302 -80 303 -79
rect 303 -80 304 -79
rect 304 -80 305 -79
rect 305 -80 306 -79
rect 306 -80 307 -79
rect 307 -80 308 -79
rect 308 -80 309 -79
rect 309 -80 310 -79
rect 310 -80 311 -79
rect 311 -80 312 -79
rect 312 -80 313 -79
rect 313 -80 314 -79
rect 314 -80 315 -79
rect 315 -80 316 -79
rect 316 -80 317 -79
rect 317 -80 318 -79
rect 318 -80 319 -79
rect 319 -80 320 -79
rect 320 -80 321 -79
rect 321 -80 322 -79
rect 322 -80 323 -79
rect 323 -80 324 -79
rect 324 -80 325 -79
rect 325 -80 326 -79
rect 326 -80 327 -79
rect 327 -80 328 -79
rect 328 -80 329 -79
rect 329 -80 330 -79
rect 330 -80 331 -79
rect 331 -80 332 -79
rect 332 -80 333 -79
rect 333 -80 334 -79
rect 334 -80 335 -79
rect 335 -80 336 -79
rect 336 -80 337 -79
rect 337 -80 338 -79
rect 338 -80 339 -79
rect 339 -80 340 -79
rect 340 -80 341 -79
rect 341 -80 342 -79
rect 342 -80 343 -79
rect 343 -80 344 -79
rect 344 -80 345 -79
rect 345 -80 346 -79
rect 346 -80 347 -79
rect 347 -80 348 -79
rect 348 -80 349 -79
rect 349 -80 350 -79
rect 350 -80 351 -79
rect 351 -80 352 -79
rect 352 -80 353 -79
rect 353 -80 354 -79
rect 354 -80 355 -79
rect 355 -80 356 -79
rect 356 -80 357 -79
rect 357 -80 358 -79
rect 358 -80 359 -79
rect 359 -80 360 -79
rect 360 -80 361 -79
rect 361 -80 362 -79
rect 362 -80 363 -79
rect 363 -80 364 -79
rect 364 -80 365 -79
rect 365 -80 366 -79
rect 366 -80 367 -79
rect 367 -80 368 -79
rect 368 -80 369 -79
rect 369 -80 370 -79
rect 370 -80 371 -79
rect 371 -80 372 -79
rect 372 -80 373 -79
rect 373 -80 374 -79
rect 374 -80 375 -79
rect 375 -80 376 -79
rect 376 -80 377 -79
rect 377 -80 378 -79
rect 378 -80 379 -79
rect 379 -80 380 -79
rect 380 -80 381 -79
rect 381 -80 382 -79
rect 382 -80 383 -79
rect 383 -80 384 -79
rect 384 -80 385 -79
rect 385 -80 386 -79
rect 386 -80 387 -79
rect 387 -80 388 -79
rect 388 -80 389 -79
rect 389 -80 390 -79
rect 390 -80 391 -79
rect 391 -80 392 -79
rect 392 -80 393 -79
rect 393 -80 394 -79
rect 394 -80 395 -79
rect 395 -80 396 -79
rect 396 -80 397 -79
rect 397 -80 398 -79
rect 398 -80 399 -79
rect 399 -80 400 -79
rect 400 -80 401 -79
rect 401 -80 402 -79
rect 402 -80 403 -79
rect 403 -80 404 -79
rect 404 -80 405 -79
rect 405 -80 406 -79
rect 406 -80 407 -79
rect 407 -80 408 -79
rect 408 -80 409 -79
rect 409 -80 410 -79
rect 410 -80 411 -79
rect 411 -80 412 -79
rect 412 -80 413 -79
rect 413 -80 414 -79
rect 414 -80 415 -79
rect 415 -80 416 -79
rect 416 -80 417 -79
rect 417 -80 418 -79
rect 418 -80 419 -79
rect 419 -80 420 -79
rect 420 -80 421 -79
rect 421 -80 422 -79
rect 422 -80 423 -79
rect 423 -80 424 -79
rect 424 -80 425 -79
rect 425 -80 426 -79
rect 426 -80 427 -79
rect 427 -80 428 -79
rect 428 -80 429 -79
rect 429 -80 430 -79
rect 430 -80 431 -79
rect 431 -80 432 -79
rect 432 -80 433 -79
rect 433 -80 434 -79
rect 434 -80 435 -79
rect 435 -80 436 -79
rect 436 -80 437 -79
rect 437 -80 438 -79
rect 438 -80 439 -79
rect 439 -80 440 -79
rect 440 -80 441 -79
rect 441 -80 442 -79
rect 442 -80 443 -79
rect 443 -80 444 -79
rect 444 -80 445 -79
rect 445 -80 446 -79
rect 446 -80 447 -79
rect 447 -80 448 -79
rect 448 -80 449 -79
rect 449 -80 450 -79
rect 450 -80 451 -79
rect 451 -80 452 -79
rect 452 -80 453 -79
rect 453 -80 454 -79
rect 454 -80 455 -79
rect 455 -80 456 -79
rect 456 -80 457 -79
rect 457 -80 458 -79
rect 458 -80 459 -79
rect 459 -80 460 -79
rect 460 -80 461 -79
rect 461 -80 462 -79
rect 462 -80 463 -79
rect 463 -80 464 -79
rect 464 -80 465 -79
rect 465 -80 466 -79
rect 466 -80 467 -79
rect 467 -80 468 -79
rect 468 -80 469 -79
rect 469 -80 470 -79
rect 470 -80 471 -79
rect 471 -80 472 -79
rect 472 -80 473 -79
rect 473 -80 474 -79
rect 474 -80 475 -79
rect 475 -80 476 -79
rect 476 -80 477 -79
rect 477 -80 478 -79
rect 478 -80 479 -79
rect 479 -80 480 -79
rect 2 -81 3 -80
rect 3 -81 4 -80
rect 4 -81 5 -80
rect 5 -81 6 -80
rect 6 -81 7 -80
rect 7 -81 8 -80
rect 8 -81 9 -80
rect 9 -81 10 -80
rect 10 -81 11 -80
rect 11 -81 12 -80
rect 12 -81 13 -80
rect 13 -81 14 -80
rect 14 -81 15 -80
rect 15 -81 16 -80
rect 16 -81 17 -80
rect 17 -81 18 -80
rect 18 -81 19 -80
rect 19 -81 20 -80
rect 20 -81 21 -80
rect 21 -81 22 -80
rect 22 -81 23 -80
rect 23 -81 24 -80
rect 24 -81 25 -80
rect 25 -81 26 -80
rect 39 -81 40 -80
rect 40 -81 41 -80
rect 41 -81 42 -80
rect 42 -81 43 -80
rect 43 -81 44 -80
rect 44 -81 45 -80
rect 45 -81 46 -80
rect 46 -81 47 -80
rect 47 -81 48 -80
rect 48 -81 49 -80
rect 49 -81 50 -80
rect 50 -81 51 -80
rect 51 -81 52 -80
rect 52 -81 53 -80
rect 53 -81 54 -80
rect 54 -81 55 -80
rect 55 -81 56 -80
rect 56 -81 57 -80
rect 57 -81 58 -80
rect 71 -81 72 -80
rect 72 -81 73 -80
rect 73 -81 74 -80
rect 74 -81 75 -80
rect 75 -81 76 -80
rect 76 -81 77 -80
rect 77 -81 78 -80
rect 78 -81 79 -80
rect 79 -81 80 -80
rect 80 -81 81 -80
rect 81 -81 82 -80
rect 82 -81 83 -80
rect 83 -81 84 -80
rect 84 -81 85 -80
rect 85 -81 86 -80
rect 86 -81 87 -80
rect 87 -81 88 -80
rect 88 -81 89 -80
rect 89 -81 90 -80
rect 103 -81 104 -80
rect 104 -81 105 -80
rect 105 -81 106 -80
rect 106 -81 107 -80
rect 107 -81 108 -80
rect 108 -81 109 -80
rect 109 -81 110 -80
rect 110 -81 111 -80
rect 111 -81 112 -80
rect 112 -81 113 -80
rect 113 -81 114 -80
rect 114 -81 115 -80
rect 115 -81 116 -80
rect 116 -81 117 -80
rect 117 -81 118 -80
rect 118 -81 119 -80
rect 119 -81 120 -80
rect 120 -81 121 -80
rect 121 -81 122 -80
rect 135 -81 136 -80
rect 136 -81 137 -80
rect 137 -81 138 -80
rect 138 -81 139 -80
rect 139 -81 140 -80
rect 140 -81 141 -80
rect 141 -81 142 -80
rect 142 -81 143 -80
rect 143 -81 144 -80
rect 144 -81 145 -80
rect 145 -81 146 -80
rect 146 -81 147 -80
rect 147 -81 148 -80
rect 148 -81 149 -80
rect 149 -81 150 -80
rect 150 -81 151 -80
rect 151 -81 152 -80
rect 152 -81 153 -80
rect 153 -81 154 -80
rect 167 -81 168 -80
rect 168 -81 169 -80
rect 169 -81 170 -80
rect 170 -81 171 -80
rect 171 -81 172 -80
rect 172 -81 173 -80
rect 173 -81 174 -80
rect 174 -81 175 -80
rect 175 -81 176 -80
rect 176 -81 177 -80
rect 177 -81 178 -80
rect 178 -81 179 -80
rect 179 -81 180 -80
rect 180 -81 181 -80
rect 181 -81 182 -80
rect 182 -81 183 -80
rect 183 -81 184 -80
rect 184 -81 185 -80
rect 185 -81 186 -80
rect 186 -81 187 -80
rect 187 -81 188 -80
rect 188 -81 189 -80
rect 189 -81 190 -80
rect 190 -81 191 -80
rect 191 -81 192 -80
rect 192 -81 193 -80
rect 193 -81 194 -80
rect 194 -81 195 -80
rect 195 -81 196 -80
rect 196 -81 197 -80
rect 197 -81 198 -80
rect 198 -81 199 -80
rect 199 -81 200 -80
rect 200 -81 201 -80
rect 201 -81 202 -80
rect 202 -81 203 -80
rect 203 -81 204 -80
rect 204 -81 205 -80
rect 205 -81 206 -80
rect 206 -81 207 -80
rect 207 -81 208 -80
rect 208 -81 209 -80
rect 209 -81 210 -80
rect 210 -81 211 -80
rect 211 -81 212 -80
rect 212 -81 213 -80
rect 213 -81 214 -80
rect 214 -81 215 -80
rect 215 -81 216 -80
rect 216 -81 217 -80
rect 217 -81 218 -80
rect 218 -81 219 -80
rect 219 -81 220 -80
rect 220 -81 221 -80
rect 221 -81 222 -80
rect 222 -81 223 -80
rect 223 -81 224 -80
rect 224 -81 225 -80
rect 225 -81 226 -80
rect 226 -81 227 -80
rect 227 -81 228 -80
rect 228 -81 229 -80
rect 229 -81 230 -80
rect 230 -81 231 -80
rect 231 -81 232 -80
rect 232 -81 233 -80
rect 233 -81 234 -80
rect 234 -81 235 -80
rect 235 -81 236 -80
rect 236 -81 237 -80
rect 237 -81 238 -80
rect 238 -81 239 -80
rect 239 -81 240 -80
rect 240 -81 241 -80
rect 241 -81 242 -80
rect 242 -81 243 -80
rect 243 -81 244 -80
rect 244 -81 245 -80
rect 245 -81 246 -80
rect 246 -81 247 -80
rect 247 -81 248 -80
rect 248 -81 249 -80
rect 249 -81 250 -80
rect 250 -81 251 -80
rect 251 -81 252 -80
rect 252 -81 253 -80
rect 253 -81 254 -80
rect 254 -81 255 -80
rect 255 -81 256 -80
rect 256 -81 257 -80
rect 257 -81 258 -80
rect 258 -81 259 -80
rect 259 -81 260 -80
rect 260 -81 261 -80
rect 261 -81 262 -80
rect 262 -81 263 -80
rect 263 -81 264 -80
rect 264 -81 265 -80
rect 265 -81 266 -80
rect 266 -81 267 -80
rect 267 -81 268 -80
rect 268 -81 269 -80
rect 269 -81 270 -80
rect 270 -81 271 -80
rect 271 -81 272 -80
rect 272 -81 273 -80
rect 273 -81 274 -80
rect 274 -81 275 -80
rect 275 -81 276 -80
rect 276 -81 277 -80
rect 277 -81 278 -80
rect 278 -81 279 -80
rect 279 -81 280 -80
rect 280 -81 281 -80
rect 281 -81 282 -80
rect 282 -81 283 -80
rect 283 -81 284 -80
rect 284 -81 285 -80
rect 285 -81 286 -80
rect 286 -81 287 -80
rect 287 -81 288 -80
rect 288 -81 289 -80
rect 289 -81 290 -80
rect 290 -81 291 -80
rect 291 -81 292 -80
rect 292 -81 293 -80
rect 293 -81 294 -80
rect 294 -81 295 -80
rect 295 -81 296 -80
rect 296 -81 297 -80
rect 297 -81 298 -80
rect 298 -81 299 -80
rect 299 -81 300 -80
rect 300 -81 301 -80
rect 301 -81 302 -80
rect 302 -81 303 -80
rect 303 -81 304 -80
rect 304 -81 305 -80
rect 305 -81 306 -80
rect 306 -81 307 -80
rect 307 -81 308 -80
rect 308 -81 309 -80
rect 309 -81 310 -80
rect 310 -81 311 -80
rect 311 -81 312 -80
rect 312 -81 313 -80
rect 313 -81 314 -80
rect 314 -81 315 -80
rect 315 -81 316 -80
rect 316 -81 317 -80
rect 317 -81 318 -80
rect 318 -81 319 -80
rect 319 -81 320 -80
rect 320 -81 321 -80
rect 321 -81 322 -80
rect 322 -81 323 -80
rect 323 -81 324 -80
rect 324 -81 325 -80
rect 325 -81 326 -80
rect 326 -81 327 -80
rect 327 -81 328 -80
rect 328 -81 329 -80
rect 329 -81 330 -80
rect 330 -81 331 -80
rect 331 -81 332 -80
rect 332 -81 333 -80
rect 333 -81 334 -80
rect 334 -81 335 -80
rect 335 -81 336 -80
rect 336 -81 337 -80
rect 337 -81 338 -80
rect 338 -81 339 -80
rect 339 -81 340 -80
rect 340 -81 341 -80
rect 341 -81 342 -80
rect 342 -81 343 -80
rect 343 -81 344 -80
rect 344 -81 345 -80
rect 345 -81 346 -80
rect 346 -81 347 -80
rect 347 -81 348 -80
rect 348 -81 349 -80
rect 349 -81 350 -80
rect 350 -81 351 -80
rect 351 -81 352 -80
rect 352 -81 353 -80
rect 353 -81 354 -80
rect 354 -81 355 -80
rect 355 -81 356 -80
rect 356 -81 357 -80
rect 357 -81 358 -80
rect 358 -81 359 -80
rect 359 -81 360 -80
rect 360 -81 361 -80
rect 361 -81 362 -80
rect 362 -81 363 -80
rect 363 -81 364 -80
rect 364 -81 365 -80
rect 365 -81 366 -80
rect 366 -81 367 -80
rect 367 -81 368 -80
rect 368 -81 369 -80
rect 369 -81 370 -80
rect 370 -81 371 -80
rect 371 -81 372 -80
rect 372 -81 373 -80
rect 373 -81 374 -80
rect 374 -81 375 -80
rect 375 -81 376 -80
rect 376 -81 377 -80
rect 377 -81 378 -80
rect 378 -81 379 -80
rect 379 -81 380 -80
rect 380 -81 381 -80
rect 381 -81 382 -80
rect 382 -81 383 -80
rect 383 -81 384 -80
rect 384 -81 385 -80
rect 385 -81 386 -80
rect 386 -81 387 -80
rect 387 -81 388 -80
rect 388 -81 389 -80
rect 389 -81 390 -80
rect 390 -81 391 -80
rect 391 -81 392 -80
rect 392 -81 393 -80
rect 393 -81 394 -80
rect 394 -81 395 -80
rect 395 -81 396 -80
rect 396 -81 397 -80
rect 397 -81 398 -80
rect 398 -81 399 -80
rect 399 -81 400 -80
rect 400 -81 401 -80
rect 401 -81 402 -80
rect 402 -81 403 -80
rect 403 -81 404 -80
rect 404 -81 405 -80
rect 405 -81 406 -80
rect 406 -81 407 -80
rect 407 -81 408 -80
rect 408 -81 409 -80
rect 409 -81 410 -80
rect 410 -81 411 -80
rect 411 -81 412 -80
rect 412 -81 413 -80
rect 413 -81 414 -80
rect 414 -81 415 -80
rect 415 -81 416 -80
rect 416 -81 417 -80
rect 417 -81 418 -80
rect 418 -81 419 -80
rect 419 -81 420 -80
rect 420 -81 421 -80
rect 421 -81 422 -80
rect 422 -81 423 -80
rect 423 -81 424 -80
rect 424 -81 425 -80
rect 425 -81 426 -80
rect 426 -81 427 -80
rect 427 -81 428 -80
rect 428 -81 429 -80
rect 429 -81 430 -80
rect 430 -81 431 -80
rect 431 -81 432 -80
rect 432 -81 433 -80
rect 433 -81 434 -80
rect 434 -81 435 -80
rect 435 -81 436 -80
rect 436 -81 437 -80
rect 437 -81 438 -80
rect 438 -81 439 -80
rect 439 -81 440 -80
rect 440 -81 441 -80
rect 441 -81 442 -80
rect 442 -81 443 -80
rect 443 -81 444 -80
rect 444 -81 445 -80
rect 445 -81 446 -80
rect 446 -81 447 -80
rect 447 -81 448 -80
rect 448 -81 449 -80
rect 449 -81 450 -80
rect 450 -81 451 -80
rect 451 -81 452 -80
rect 452 -81 453 -80
rect 453 -81 454 -80
rect 454 -81 455 -80
rect 455 -81 456 -80
rect 456 -81 457 -80
rect 457 -81 458 -80
rect 458 -81 459 -80
rect 459 -81 460 -80
rect 460 -81 461 -80
rect 461 -81 462 -80
rect 462 -81 463 -80
rect 463 -81 464 -80
rect 464 -81 465 -80
rect 465 -81 466 -80
rect 466 -81 467 -80
rect 467 -81 468 -80
rect 468 -81 469 -80
rect 469 -81 470 -80
rect 470 -81 471 -80
rect 471 -81 472 -80
rect 472 -81 473 -80
rect 473 -81 474 -80
rect 474 -81 475 -80
rect 475 -81 476 -80
rect 476 -81 477 -80
rect 477 -81 478 -80
rect 478 -81 479 -80
rect 479 -81 480 -80
rect 2 -82 3 -81
rect 3 -82 4 -81
rect 4 -82 5 -81
rect 5 -82 6 -81
rect 6 -82 7 -81
rect 7 -82 8 -81
rect 8 -82 9 -81
rect 9 -82 10 -81
rect 10 -82 11 -81
rect 11 -82 12 -81
rect 12 -82 13 -81
rect 13 -82 14 -81
rect 14 -82 15 -81
rect 15 -82 16 -81
rect 16 -82 17 -81
rect 17 -82 18 -81
rect 18 -82 19 -81
rect 19 -82 20 -81
rect 20 -82 21 -81
rect 21 -82 22 -81
rect 22 -82 23 -81
rect 23 -82 24 -81
rect 24 -82 25 -81
rect 25 -82 26 -81
rect 26 -82 27 -81
rect 27 -82 28 -81
rect 38 -82 39 -81
rect 39 -82 40 -81
rect 40 -82 41 -81
rect 41 -82 42 -81
rect 42 -82 43 -81
rect 43 -82 44 -81
rect 44 -82 45 -81
rect 45 -82 46 -81
rect 46 -82 47 -81
rect 47 -82 48 -81
rect 48 -82 49 -81
rect 49 -82 50 -81
rect 50 -82 51 -81
rect 51 -82 52 -81
rect 52 -82 53 -81
rect 53 -82 54 -81
rect 54 -82 55 -81
rect 55 -82 56 -81
rect 56 -82 57 -81
rect 57 -82 58 -81
rect 58 -82 59 -81
rect 59 -82 60 -81
rect 70 -82 71 -81
rect 71 -82 72 -81
rect 72 -82 73 -81
rect 73 -82 74 -81
rect 74 -82 75 -81
rect 75 -82 76 -81
rect 76 -82 77 -81
rect 77 -82 78 -81
rect 78 -82 79 -81
rect 79 -82 80 -81
rect 80 -82 81 -81
rect 81 -82 82 -81
rect 82 -82 83 -81
rect 83 -82 84 -81
rect 84 -82 85 -81
rect 85 -82 86 -81
rect 86 -82 87 -81
rect 87 -82 88 -81
rect 88 -82 89 -81
rect 89 -82 90 -81
rect 90 -82 91 -81
rect 91 -82 92 -81
rect 102 -82 103 -81
rect 103 -82 104 -81
rect 104 -82 105 -81
rect 105 -82 106 -81
rect 106 -82 107 -81
rect 107 -82 108 -81
rect 108 -82 109 -81
rect 109 -82 110 -81
rect 110 -82 111 -81
rect 111 -82 112 -81
rect 112 -82 113 -81
rect 113 -82 114 -81
rect 114 -82 115 -81
rect 115 -82 116 -81
rect 116 -82 117 -81
rect 117 -82 118 -81
rect 118 -82 119 -81
rect 119 -82 120 -81
rect 120 -82 121 -81
rect 121 -82 122 -81
rect 122 -82 123 -81
rect 123 -82 124 -81
rect 134 -82 135 -81
rect 135 -82 136 -81
rect 136 -82 137 -81
rect 137 -82 138 -81
rect 138 -82 139 -81
rect 139 -82 140 -81
rect 140 -82 141 -81
rect 141 -82 142 -81
rect 142 -82 143 -81
rect 143 -82 144 -81
rect 144 -82 145 -81
rect 145 -82 146 -81
rect 146 -82 147 -81
rect 147 -82 148 -81
rect 148 -82 149 -81
rect 149 -82 150 -81
rect 150 -82 151 -81
rect 151 -82 152 -81
rect 152 -82 153 -81
rect 153 -82 154 -81
rect 154 -82 155 -81
rect 155 -82 156 -81
rect 166 -82 167 -81
rect 167 -82 168 -81
rect 168 -82 169 -81
rect 169 -82 170 -81
rect 170 -82 171 -81
rect 171 -82 172 -81
rect 172 -82 173 -81
rect 173 -82 174 -81
rect 174 -82 175 -81
rect 175 -82 176 -81
rect 176 -82 177 -81
rect 177 -82 178 -81
rect 178 -82 179 -81
rect 179 -82 180 -81
rect 180 -82 181 -81
rect 181 -82 182 -81
rect 182 -82 183 -81
rect 183 -82 184 -81
rect 184 -82 185 -81
rect 185 -82 186 -81
rect 186 -82 187 -81
rect 187 -82 188 -81
rect 188 -82 189 -81
rect 189 -82 190 -81
rect 190 -82 191 -81
rect 191 -82 192 -81
rect 192 -82 193 -81
rect 193 -82 194 -81
rect 194 -82 195 -81
rect 195 -82 196 -81
rect 196 -82 197 -81
rect 197 -82 198 -81
rect 198 -82 199 -81
rect 199 -82 200 -81
rect 200 -82 201 -81
rect 201 -82 202 -81
rect 202 -82 203 -81
rect 203 -82 204 -81
rect 204 -82 205 -81
rect 205 -82 206 -81
rect 206 -82 207 -81
rect 207 -82 208 -81
rect 208 -82 209 -81
rect 209 -82 210 -81
rect 210 -82 211 -81
rect 211 -82 212 -81
rect 212 -82 213 -81
rect 213 -82 214 -81
rect 214 -82 215 -81
rect 215 -82 216 -81
rect 216 -82 217 -81
rect 217 -82 218 -81
rect 218 -82 219 -81
rect 219 -82 220 -81
rect 220 -82 221 -81
rect 221 -82 222 -81
rect 222 -82 223 -81
rect 223 -82 224 -81
rect 224 -82 225 -81
rect 225 -82 226 -81
rect 226 -82 227 -81
rect 227 -82 228 -81
rect 228 -82 229 -81
rect 229 -82 230 -81
rect 230 -82 231 -81
rect 231 -82 232 -81
rect 232 -82 233 -81
rect 233 -82 234 -81
rect 234 -82 235 -81
rect 235 -82 236 -81
rect 236 -82 237 -81
rect 237 -82 238 -81
rect 238 -82 239 -81
rect 239 -82 240 -81
rect 240 -82 241 -81
rect 241 -82 242 -81
rect 242 -82 243 -81
rect 243 -82 244 -81
rect 244 -82 245 -81
rect 245 -82 246 -81
rect 246 -82 247 -81
rect 247 -82 248 -81
rect 248 -82 249 -81
rect 249 -82 250 -81
rect 250 -82 251 -81
rect 251 -82 252 -81
rect 252 -82 253 -81
rect 253 -82 254 -81
rect 254 -82 255 -81
rect 255 -82 256 -81
rect 256 -82 257 -81
rect 257 -82 258 -81
rect 258 -82 259 -81
rect 259 -82 260 -81
rect 260 -82 261 -81
rect 261 -82 262 -81
rect 262 -82 263 -81
rect 263 -82 264 -81
rect 264 -82 265 -81
rect 265 -82 266 -81
rect 266 -82 267 -81
rect 267 -82 268 -81
rect 268 -82 269 -81
rect 269 -82 270 -81
rect 270 -82 271 -81
rect 271 -82 272 -81
rect 272 -82 273 -81
rect 273 -82 274 -81
rect 274 -82 275 -81
rect 275 -82 276 -81
rect 276 -82 277 -81
rect 277 -82 278 -81
rect 278 -82 279 -81
rect 279 -82 280 -81
rect 280 -82 281 -81
rect 281 -82 282 -81
rect 282 -82 283 -81
rect 283 -82 284 -81
rect 284 -82 285 -81
rect 285 -82 286 -81
rect 286 -82 287 -81
rect 287 -82 288 -81
rect 288 -82 289 -81
rect 289 -82 290 -81
rect 290 -82 291 -81
rect 291 -82 292 -81
rect 292 -82 293 -81
rect 293 -82 294 -81
rect 294 -82 295 -81
rect 295 -82 296 -81
rect 296 -82 297 -81
rect 297 -82 298 -81
rect 298 -82 299 -81
rect 299 -82 300 -81
rect 300 -82 301 -81
rect 301 -82 302 -81
rect 302 -82 303 -81
rect 303 -82 304 -81
rect 304 -82 305 -81
rect 305 -82 306 -81
rect 306 -82 307 -81
rect 307 -82 308 -81
rect 308 -82 309 -81
rect 309 -82 310 -81
rect 310 -82 311 -81
rect 311 -82 312 -81
rect 312 -82 313 -81
rect 313 -82 314 -81
rect 314 -82 315 -81
rect 315 -82 316 -81
rect 316 -82 317 -81
rect 317 -82 318 -81
rect 318 -82 319 -81
rect 319 -82 320 -81
rect 320 -82 321 -81
rect 321 -82 322 -81
rect 322 -82 323 -81
rect 323 -82 324 -81
rect 324 -82 325 -81
rect 325 -82 326 -81
rect 326 -82 327 -81
rect 327 -82 328 -81
rect 328 -82 329 -81
rect 329 -82 330 -81
rect 330 -82 331 -81
rect 331 -82 332 -81
rect 332 -82 333 -81
rect 333 -82 334 -81
rect 334 -82 335 -81
rect 335 -82 336 -81
rect 336 -82 337 -81
rect 337 -82 338 -81
rect 338 -82 339 -81
rect 339 -82 340 -81
rect 340 -82 341 -81
rect 341 -82 342 -81
rect 342 -82 343 -81
rect 343 -82 344 -81
rect 344 -82 345 -81
rect 345 -82 346 -81
rect 346 -82 347 -81
rect 347 -82 348 -81
rect 348 -82 349 -81
rect 349 -82 350 -81
rect 350 -82 351 -81
rect 351 -82 352 -81
rect 352 -82 353 -81
rect 353 -82 354 -81
rect 354 -82 355 -81
rect 355 -82 356 -81
rect 356 -82 357 -81
rect 357 -82 358 -81
rect 358 -82 359 -81
rect 359 -82 360 -81
rect 360 -82 361 -81
rect 361 -82 362 -81
rect 362 -82 363 -81
rect 363 -82 364 -81
rect 364 -82 365 -81
rect 365 -82 366 -81
rect 366 -82 367 -81
rect 367 -82 368 -81
rect 368 -82 369 -81
rect 369 -82 370 -81
rect 370 -82 371 -81
rect 371 -82 372 -81
rect 372 -82 373 -81
rect 373 -82 374 -81
rect 374 -82 375 -81
rect 375 -82 376 -81
rect 376 -82 377 -81
rect 377 -82 378 -81
rect 378 -82 379 -81
rect 379 -82 380 -81
rect 380 -82 381 -81
rect 381 -82 382 -81
rect 382 -82 383 -81
rect 383 -82 384 -81
rect 384 -82 385 -81
rect 385 -82 386 -81
rect 386 -82 387 -81
rect 387 -82 388 -81
rect 388 -82 389 -81
rect 389 -82 390 -81
rect 390 -82 391 -81
rect 391 -82 392 -81
rect 392 -82 393 -81
rect 393 -82 394 -81
rect 394 -82 395 -81
rect 395 -82 396 -81
rect 396 -82 397 -81
rect 397 -82 398 -81
rect 398 -82 399 -81
rect 399 -82 400 -81
rect 400 -82 401 -81
rect 401 -82 402 -81
rect 402 -82 403 -81
rect 403 -82 404 -81
rect 404 -82 405 -81
rect 405 -82 406 -81
rect 406 -82 407 -81
rect 407 -82 408 -81
rect 408 -82 409 -81
rect 409 -82 410 -81
rect 410 -82 411 -81
rect 411 -82 412 -81
rect 412 -82 413 -81
rect 413 -82 414 -81
rect 414 -82 415 -81
rect 415 -82 416 -81
rect 416 -82 417 -81
rect 417 -82 418 -81
rect 418 -82 419 -81
rect 419 -82 420 -81
rect 420 -82 421 -81
rect 421 -82 422 -81
rect 422 -82 423 -81
rect 423 -82 424 -81
rect 424 -82 425 -81
rect 425 -82 426 -81
rect 426 -82 427 -81
rect 427 -82 428 -81
rect 428 -82 429 -81
rect 429 -82 430 -81
rect 430 -82 431 -81
rect 431 -82 432 -81
rect 432 -82 433 -81
rect 433 -82 434 -81
rect 434 -82 435 -81
rect 435 -82 436 -81
rect 436 -82 437 -81
rect 437 -82 438 -81
rect 438 -82 439 -81
rect 439 -82 440 -81
rect 440 -82 441 -81
rect 441 -82 442 -81
rect 442 -82 443 -81
rect 443 -82 444 -81
rect 444 -82 445 -81
rect 445 -82 446 -81
rect 446 -82 447 -81
rect 447 -82 448 -81
rect 448 -82 449 -81
rect 449 -82 450 -81
rect 450 -82 451 -81
rect 451 -82 452 -81
rect 452 -82 453 -81
rect 453 -82 454 -81
rect 454 -82 455 -81
rect 455 -82 456 -81
rect 456 -82 457 -81
rect 457 -82 458 -81
rect 458 -82 459 -81
rect 459 -82 460 -81
rect 460 -82 461 -81
rect 461 -82 462 -81
rect 462 -82 463 -81
rect 463 -82 464 -81
rect 464 -82 465 -81
rect 465 -82 466 -81
rect 466 -82 467 -81
rect 467 -82 468 -81
rect 468 -82 469 -81
rect 469 -82 470 -81
rect 470 -82 471 -81
rect 471 -82 472 -81
rect 472 -82 473 -81
rect 473 -82 474 -81
rect 474 -82 475 -81
rect 475 -82 476 -81
rect 476 -82 477 -81
rect 477 -82 478 -81
rect 478 -82 479 -81
rect 479 -82 480 -81
rect 2 -83 3 -82
rect 3 -83 4 -82
rect 4 -83 5 -82
rect 5 -83 6 -82
rect 6 -83 7 -82
rect 7 -83 8 -82
rect 8 -83 9 -82
rect 9 -83 10 -82
rect 10 -83 11 -82
rect 11 -83 12 -82
rect 12 -83 13 -82
rect 13 -83 14 -82
rect 14 -83 15 -82
rect 15 -83 16 -82
rect 16 -83 17 -82
rect 17 -83 18 -82
rect 18 -83 19 -82
rect 19 -83 20 -82
rect 20 -83 21 -82
rect 21 -83 22 -82
rect 22 -83 23 -82
rect 23 -83 24 -82
rect 24 -83 25 -82
rect 25 -83 26 -82
rect 26 -83 27 -82
rect 27 -83 28 -82
rect 37 -83 38 -82
rect 38 -83 39 -82
rect 39 -83 40 -82
rect 40 -83 41 -82
rect 41 -83 42 -82
rect 42 -83 43 -82
rect 43 -83 44 -82
rect 44 -83 45 -82
rect 45 -83 46 -82
rect 46 -83 47 -82
rect 47 -83 48 -82
rect 48 -83 49 -82
rect 49 -83 50 -82
rect 50 -83 51 -82
rect 51 -83 52 -82
rect 52 -83 53 -82
rect 53 -83 54 -82
rect 54 -83 55 -82
rect 55 -83 56 -82
rect 56 -83 57 -82
rect 57 -83 58 -82
rect 58 -83 59 -82
rect 59 -83 60 -82
rect 69 -83 70 -82
rect 70 -83 71 -82
rect 71 -83 72 -82
rect 72 -83 73 -82
rect 73 -83 74 -82
rect 74 -83 75 -82
rect 75 -83 76 -82
rect 76 -83 77 -82
rect 77 -83 78 -82
rect 78 -83 79 -82
rect 79 -83 80 -82
rect 80 -83 81 -82
rect 81 -83 82 -82
rect 82 -83 83 -82
rect 83 -83 84 -82
rect 84 -83 85 -82
rect 85 -83 86 -82
rect 86 -83 87 -82
rect 87 -83 88 -82
rect 88 -83 89 -82
rect 89 -83 90 -82
rect 90 -83 91 -82
rect 91 -83 92 -82
rect 101 -83 102 -82
rect 102 -83 103 -82
rect 103 -83 104 -82
rect 104 -83 105 -82
rect 105 -83 106 -82
rect 106 -83 107 -82
rect 107 -83 108 -82
rect 108 -83 109 -82
rect 109 -83 110 -82
rect 110 -83 111 -82
rect 111 -83 112 -82
rect 112 -83 113 -82
rect 113 -83 114 -82
rect 114 -83 115 -82
rect 115 -83 116 -82
rect 116 -83 117 -82
rect 117 -83 118 -82
rect 118 -83 119 -82
rect 119 -83 120 -82
rect 120 -83 121 -82
rect 121 -83 122 -82
rect 122 -83 123 -82
rect 123 -83 124 -82
rect 133 -83 134 -82
rect 134 -83 135 -82
rect 135 -83 136 -82
rect 136 -83 137 -82
rect 137 -83 138 -82
rect 138 -83 139 -82
rect 139 -83 140 -82
rect 140 -83 141 -82
rect 141 -83 142 -82
rect 142 -83 143 -82
rect 143 -83 144 -82
rect 144 -83 145 -82
rect 145 -83 146 -82
rect 146 -83 147 -82
rect 147 -83 148 -82
rect 148 -83 149 -82
rect 149 -83 150 -82
rect 150 -83 151 -82
rect 151 -83 152 -82
rect 152 -83 153 -82
rect 153 -83 154 -82
rect 154 -83 155 -82
rect 155 -83 156 -82
rect 165 -83 166 -82
rect 166 -83 167 -82
rect 167 -83 168 -82
rect 168 -83 169 -82
rect 169 -83 170 -82
rect 170 -83 171 -82
rect 171 -83 172 -82
rect 172 -83 173 -82
rect 173 -83 174 -82
rect 174 -83 175 -82
rect 175 -83 176 -82
rect 176 -83 177 -82
rect 177 -83 178 -82
rect 178 -83 179 -82
rect 179 -83 180 -82
rect 180 -83 181 -82
rect 181 -83 182 -82
rect 182 -83 183 -82
rect 183 -83 184 -82
rect 184 -83 185 -82
rect 185 -83 186 -82
rect 186 -83 187 -82
rect 187 -83 188 -82
rect 188 -83 189 -82
rect 189 -83 190 -82
rect 190 -83 191 -82
rect 191 -83 192 -82
rect 192 -83 193 -82
rect 193 -83 194 -82
rect 194 -83 195 -82
rect 195 -83 196 -82
rect 196 -83 197 -82
rect 197 -83 198 -82
rect 198 -83 199 -82
rect 199 -83 200 -82
rect 200 -83 201 -82
rect 201 -83 202 -82
rect 202 -83 203 -82
rect 203 -83 204 -82
rect 204 -83 205 -82
rect 205 -83 206 -82
rect 206 -83 207 -82
rect 207 -83 208 -82
rect 208 -83 209 -82
rect 209 -83 210 -82
rect 210 -83 211 -82
rect 211 -83 212 -82
rect 212 -83 213 -82
rect 213 -83 214 -82
rect 214 -83 215 -82
rect 215 -83 216 -82
rect 216 -83 217 -82
rect 217 -83 218 -82
rect 218 -83 219 -82
rect 219 -83 220 -82
rect 220 -83 221 -82
rect 221 -83 222 -82
rect 222 -83 223 -82
rect 223 -83 224 -82
rect 224 -83 225 -82
rect 225 -83 226 -82
rect 226 -83 227 -82
rect 227 -83 228 -82
rect 228 -83 229 -82
rect 229 -83 230 -82
rect 230 -83 231 -82
rect 231 -83 232 -82
rect 232 -83 233 -82
rect 233 -83 234 -82
rect 234 -83 235 -82
rect 235 -83 236 -82
rect 236 -83 237 -82
rect 237 -83 238 -82
rect 238 -83 239 -82
rect 239 -83 240 -82
rect 240 -83 241 -82
rect 241 -83 242 -82
rect 242 -83 243 -82
rect 243 -83 244 -82
rect 244 -83 245 -82
rect 245 -83 246 -82
rect 246 -83 247 -82
rect 247 -83 248 -82
rect 248 -83 249 -82
rect 249 -83 250 -82
rect 250 -83 251 -82
rect 251 -83 252 -82
rect 252 -83 253 -82
rect 253 -83 254 -82
rect 254 -83 255 -82
rect 255 -83 256 -82
rect 256 -83 257 -82
rect 257 -83 258 -82
rect 258 -83 259 -82
rect 259 -83 260 -82
rect 260 -83 261 -82
rect 261 -83 262 -82
rect 262 -83 263 -82
rect 263 -83 264 -82
rect 264 -83 265 -82
rect 265 -83 266 -82
rect 266 -83 267 -82
rect 267 -83 268 -82
rect 268 -83 269 -82
rect 269 -83 270 -82
rect 270 -83 271 -82
rect 271 -83 272 -82
rect 272 -83 273 -82
rect 273 -83 274 -82
rect 274 -83 275 -82
rect 275 -83 276 -82
rect 276 -83 277 -82
rect 277 -83 278 -82
rect 278 -83 279 -82
rect 279 -83 280 -82
rect 280 -83 281 -82
rect 281 -83 282 -82
rect 282 -83 283 -82
rect 283 -83 284 -82
rect 284 -83 285 -82
rect 285 -83 286 -82
rect 286 -83 287 -82
rect 287 -83 288 -82
rect 288 -83 289 -82
rect 289 -83 290 -82
rect 290 -83 291 -82
rect 291 -83 292 -82
rect 292 -83 293 -82
rect 293 -83 294 -82
rect 294 -83 295 -82
rect 295 -83 296 -82
rect 296 -83 297 -82
rect 297 -83 298 -82
rect 298 -83 299 -82
rect 299 -83 300 -82
rect 300 -83 301 -82
rect 301 -83 302 -82
rect 302 -83 303 -82
rect 303 -83 304 -82
rect 304 -83 305 -82
rect 305 -83 306 -82
rect 306 -83 307 -82
rect 307 -83 308 -82
rect 308 -83 309 -82
rect 309 -83 310 -82
rect 310 -83 311 -82
rect 311 -83 312 -82
rect 312 -83 313 -82
rect 313 -83 314 -82
rect 314 -83 315 -82
rect 315 -83 316 -82
rect 316 -83 317 -82
rect 317 -83 318 -82
rect 318 -83 319 -82
rect 319 -83 320 -82
rect 320 -83 321 -82
rect 321 -83 322 -82
rect 322 -83 323 -82
rect 323 -83 324 -82
rect 324 -83 325 -82
rect 325 -83 326 -82
rect 326 -83 327 -82
rect 327 -83 328 -82
rect 328 -83 329 -82
rect 329 -83 330 -82
rect 330 -83 331 -82
rect 331 -83 332 -82
rect 332 -83 333 -82
rect 333 -83 334 -82
rect 334 -83 335 -82
rect 335 -83 336 -82
rect 336 -83 337 -82
rect 337 -83 338 -82
rect 338 -83 339 -82
rect 339 -83 340 -82
rect 340 -83 341 -82
rect 341 -83 342 -82
rect 342 -83 343 -82
rect 343 -83 344 -82
rect 344 -83 345 -82
rect 345 -83 346 -82
rect 346 -83 347 -82
rect 347 -83 348 -82
rect 348 -83 349 -82
rect 349 -83 350 -82
rect 350 -83 351 -82
rect 351 -83 352 -82
rect 352 -83 353 -82
rect 353 -83 354 -82
rect 354 -83 355 -82
rect 355 -83 356 -82
rect 356 -83 357 -82
rect 357 -83 358 -82
rect 358 -83 359 -82
rect 359 -83 360 -82
rect 360 -83 361 -82
rect 361 -83 362 -82
rect 362 -83 363 -82
rect 363 -83 364 -82
rect 364 -83 365 -82
rect 365 -83 366 -82
rect 366 -83 367 -82
rect 367 -83 368 -82
rect 368 -83 369 -82
rect 369 -83 370 -82
rect 370 -83 371 -82
rect 371 -83 372 -82
rect 372 -83 373 -82
rect 373 -83 374 -82
rect 374 -83 375 -82
rect 375 -83 376 -82
rect 376 -83 377 -82
rect 377 -83 378 -82
rect 378 -83 379 -82
rect 379 -83 380 -82
rect 380 -83 381 -82
rect 381 -83 382 -82
rect 382 -83 383 -82
rect 383 -83 384 -82
rect 384 -83 385 -82
rect 385 -83 386 -82
rect 386 -83 387 -82
rect 387 -83 388 -82
rect 388 -83 389 -82
rect 389 -83 390 -82
rect 390 -83 391 -82
rect 391 -83 392 -82
rect 392 -83 393 -82
rect 393 -83 394 -82
rect 394 -83 395 -82
rect 395 -83 396 -82
rect 396 -83 397 -82
rect 397 -83 398 -82
rect 398 -83 399 -82
rect 399 -83 400 -82
rect 400 -83 401 -82
rect 401 -83 402 -82
rect 402 -83 403 -82
rect 403 -83 404 -82
rect 404 -83 405 -82
rect 405 -83 406 -82
rect 406 -83 407 -82
rect 407 -83 408 -82
rect 408 -83 409 -82
rect 409 -83 410 -82
rect 410 -83 411 -82
rect 411 -83 412 -82
rect 412 -83 413 -82
rect 413 -83 414 -82
rect 414 -83 415 -82
rect 415 -83 416 -82
rect 416 -83 417 -82
rect 417 -83 418 -82
rect 418 -83 419 -82
rect 419 -83 420 -82
rect 420 -83 421 -82
rect 421 -83 422 -82
rect 422 -83 423 -82
rect 423 -83 424 -82
rect 424 -83 425 -82
rect 425 -83 426 -82
rect 426 -83 427 -82
rect 427 -83 428 -82
rect 428 -83 429 -82
rect 429 -83 430 -82
rect 430 -83 431 -82
rect 431 -83 432 -82
rect 432 -83 433 -82
rect 433 -83 434 -82
rect 434 -83 435 -82
rect 435 -83 436 -82
rect 436 -83 437 -82
rect 437 -83 438 -82
rect 438 -83 439 -82
rect 439 -83 440 -82
rect 440 -83 441 -82
rect 441 -83 442 -82
rect 442 -83 443 -82
rect 443 -83 444 -82
rect 444 -83 445 -82
rect 445 -83 446 -82
rect 446 -83 447 -82
rect 447 -83 448 -82
rect 448 -83 449 -82
rect 449 -83 450 -82
rect 450 -83 451 -82
rect 451 -83 452 -82
rect 452 -83 453 -82
rect 453 -83 454 -82
rect 454 -83 455 -82
rect 455 -83 456 -82
rect 456 -83 457 -82
rect 457 -83 458 -82
rect 458 -83 459 -82
rect 459 -83 460 -82
rect 460 -83 461 -82
rect 461 -83 462 -82
rect 462 -83 463 -82
rect 463 -83 464 -82
rect 464 -83 465 -82
rect 465 -83 466 -82
rect 466 -83 467 -82
rect 467 -83 468 -82
rect 468 -83 469 -82
rect 469 -83 470 -82
rect 470 -83 471 -82
rect 471 -83 472 -82
rect 472 -83 473 -82
rect 473 -83 474 -82
rect 474 -83 475 -82
rect 475 -83 476 -82
rect 476 -83 477 -82
rect 477 -83 478 -82
rect 478 -83 479 -82
rect 479 -83 480 -82
rect 2 -84 3 -83
rect 3 -84 4 -83
rect 4 -84 5 -83
rect 5 -84 6 -83
rect 6 -84 7 -83
rect 7 -84 8 -83
rect 8 -84 9 -83
rect 9 -84 10 -83
rect 10 -84 11 -83
rect 11 -84 12 -83
rect 12 -84 13 -83
rect 13 -84 14 -83
rect 14 -84 15 -83
rect 15 -84 16 -83
rect 16 -84 17 -83
rect 17 -84 18 -83
rect 18 -84 19 -83
rect 19 -84 20 -83
rect 20 -84 21 -83
rect 21 -84 22 -83
rect 22 -84 23 -83
rect 23 -84 24 -83
rect 24 -84 25 -83
rect 25 -84 26 -83
rect 26 -84 27 -83
rect 27 -84 28 -83
rect 37 -84 38 -83
rect 38 -84 39 -83
rect 39 -84 40 -83
rect 40 -84 41 -83
rect 41 -84 42 -83
rect 42 -84 43 -83
rect 43 -84 44 -83
rect 44 -84 45 -83
rect 45 -84 46 -83
rect 46 -84 47 -83
rect 47 -84 48 -83
rect 48 -84 49 -83
rect 49 -84 50 -83
rect 50 -84 51 -83
rect 51 -84 52 -83
rect 52 -84 53 -83
rect 53 -84 54 -83
rect 54 -84 55 -83
rect 55 -84 56 -83
rect 56 -84 57 -83
rect 57 -84 58 -83
rect 58 -84 59 -83
rect 59 -84 60 -83
rect 69 -84 70 -83
rect 70 -84 71 -83
rect 71 -84 72 -83
rect 72 -84 73 -83
rect 73 -84 74 -83
rect 74 -84 75 -83
rect 75 -84 76 -83
rect 76 -84 77 -83
rect 77 -84 78 -83
rect 78 -84 79 -83
rect 79 -84 80 -83
rect 80 -84 81 -83
rect 81 -84 82 -83
rect 82 -84 83 -83
rect 83 -84 84 -83
rect 84 -84 85 -83
rect 85 -84 86 -83
rect 86 -84 87 -83
rect 87 -84 88 -83
rect 88 -84 89 -83
rect 89 -84 90 -83
rect 90 -84 91 -83
rect 91 -84 92 -83
rect 101 -84 102 -83
rect 102 -84 103 -83
rect 103 -84 104 -83
rect 104 -84 105 -83
rect 105 -84 106 -83
rect 106 -84 107 -83
rect 107 -84 108 -83
rect 108 -84 109 -83
rect 109 -84 110 -83
rect 110 -84 111 -83
rect 111 -84 112 -83
rect 112 -84 113 -83
rect 113 -84 114 -83
rect 114 -84 115 -83
rect 115 -84 116 -83
rect 116 -84 117 -83
rect 117 -84 118 -83
rect 118 -84 119 -83
rect 119 -84 120 -83
rect 120 -84 121 -83
rect 121 -84 122 -83
rect 122 -84 123 -83
rect 123 -84 124 -83
rect 133 -84 134 -83
rect 134 -84 135 -83
rect 135 -84 136 -83
rect 136 -84 137 -83
rect 137 -84 138 -83
rect 138 -84 139 -83
rect 139 -84 140 -83
rect 140 -84 141 -83
rect 141 -84 142 -83
rect 142 -84 143 -83
rect 143 -84 144 -83
rect 144 -84 145 -83
rect 145 -84 146 -83
rect 146 -84 147 -83
rect 147 -84 148 -83
rect 148 -84 149 -83
rect 149 -84 150 -83
rect 150 -84 151 -83
rect 151 -84 152 -83
rect 152 -84 153 -83
rect 153 -84 154 -83
rect 154 -84 155 -83
rect 155 -84 156 -83
rect 165 -84 166 -83
rect 166 -84 167 -83
rect 167 -84 168 -83
rect 168 -84 169 -83
rect 169 -84 170 -83
rect 170 -84 171 -83
rect 171 -84 172 -83
rect 172 -84 173 -83
rect 173 -84 174 -83
rect 174 -84 175 -83
rect 175 -84 176 -83
rect 176 -84 177 -83
rect 177 -84 178 -83
rect 178 -84 179 -83
rect 179 -84 180 -83
rect 180 -84 181 -83
rect 181 -84 182 -83
rect 182 -84 183 -83
rect 183 -84 184 -83
rect 184 -84 185 -83
rect 185 -84 186 -83
rect 186 -84 187 -83
rect 187 -84 188 -83
rect 188 -84 189 -83
rect 189 -84 190 -83
rect 190 -84 191 -83
rect 191 -84 192 -83
rect 192 -84 193 -83
rect 193 -84 194 -83
rect 194 -84 195 -83
rect 195 -84 196 -83
rect 196 -84 197 -83
rect 197 -84 198 -83
rect 198 -84 199 -83
rect 199 -84 200 -83
rect 200 -84 201 -83
rect 201 -84 202 -83
rect 202 -84 203 -83
rect 203 -84 204 -83
rect 204 -84 205 -83
rect 205 -84 206 -83
rect 206 -84 207 -83
rect 207 -84 208 -83
rect 208 -84 209 -83
rect 209 -84 210 -83
rect 210 -84 211 -83
rect 211 -84 212 -83
rect 212 -84 213 -83
rect 213 -84 214 -83
rect 214 -84 215 -83
rect 215 -84 216 -83
rect 216 -84 217 -83
rect 217 -84 218 -83
rect 218 -84 219 -83
rect 219 -84 220 -83
rect 220 -84 221 -83
rect 221 -84 222 -83
rect 222 -84 223 -83
rect 223 -84 224 -83
rect 224 -84 225 -83
rect 225 -84 226 -83
rect 226 -84 227 -83
rect 227 -84 228 -83
rect 228 -84 229 -83
rect 229 -84 230 -83
rect 230 -84 231 -83
rect 231 -84 232 -83
rect 232 -84 233 -83
rect 233 -84 234 -83
rect 234 -84 235 -83
rect 235 -84 236 -83
rect 236 -84 237 -83
rect 237 -84 238 -83
rect 238 -84 239 -83
rect 239 -84 240 -83
rect 240 -84 241 -83
rect 241 -84 242 -83
rect 242 -84 243 -83
rect 243 -84 244 -83
rect 244 -84 245 -83
rect 245 -84 246 -83
rect 246 -84 247 -83
rect 247 -84 248 -83
rect 248 -84 249 -83
rect 249 -84 250 -83
rect 250 -84 251 -83
rect 251 -84 252 -83
rect 252 -84 253 -83
rect 253 -84 254 -83
rect 254 -84 255 -83
rect 255 -84 256 -83
rect 256 -84 257 -83
rect 257 -84 258 -83
rect 258 -84 259 -83
rect 259 -84 260 -83
rect 260 -84 261 -83
rect 261 -84 262 -83
rect 262 -84 263 -83
rect 263 -84 264 -83
rect 264 -84 265 -83
rect 265 -84 266 -83
rect 266 -84 267 -83
rect 267 -84 268 -83
rect 268 -84 269 -83
rect 269 -84 270 -83
rect 270 -84 271 -83
rect 271 -84 272 -83
rect 272 -84 273 -83
rect 273 -84 274 -83
rect 274 -84 275 -83
rect 275 -84 276 -83
rect 276 -84 277 -83
rect 277 -84 278 -83
rect 278 -84 279 -83
rect 279 -84 280 -83
rect 280 -84 281 -83
rect 281 -84 282 -83
rect 282 -84 283 -83
rect 283 -84 284 -83
rect 284 -84 285 -83
rect 285 -84 286 -83
rect 286 -84 287 -83
rect 287 -84 288 -83
rect 288 -84 289 -83
rect 289 -84 290 -83
rect 290 -84 291 -83
rect 291 -84 292 -83
rect 292 -84 293 -83
rect 293 -84 294 -83
rect 294 -84 295 -83
rect 295 -84 296 -83
rect 296 -84 297 -83
rect 297 -84 298 -83
rect 298 -84 299 -83
rect 299 -84 300 -83
rect 300 -84 301 -83
rect 301 -84 302 -83
rect 302 -84 303 -83
rect 303 -84 304 -83
rect 304 -84 305 -83
rect 305 -84 306 -83
rect 306 -84 307 -83
rect 307 -84 308 -83
rect 308 -84 309 -83
rect 309 -84 310 -83
rect 310 -84 311 -83
rect 311 -84 312 -83
rect 312 -84 313 -83
rect 313 -84 314 -83
rect 314 -84 315 -83
rect 315 -84 316 -83
rect 316 -84 317 -83
rect 317 -84 318 -83
rect 318 -84 319 -83
rect 319 -84 320 -83
rect 320 -84 321 -83
rect 321 -84 322 -83
rect 322 -84 323 -83
rect 323 -84 324 -83
rect 324 -84 325 -83
rect 325 -84 326 -83
rect 326 -84 327 -83
rect 327 -84 328 -83
rect 328 -84 329 -83
rect 329 -84 330 -83
rect 330 -84 331 -83
rect 331 -84 332 -83
rect 332 -84 333 -83
rect 333 -84 334 -83
rect 334 -84 335 -83
rect 335 -84 336 -83
rect 336 -84 337 -83
rect 337 -84 338 -83
rect 338 -84 339 -83
rect 339 -84 340 -83
rect 340 -84 341 -83
rect 341 -84 342 -83
rect 342 -84 343 -83
rect 343 -84 344 -83
rect 344 -84 345 -83
rect 345 -84 346 -83
rect 346 -84 347 -83
rect 347 -84 348 -83
rect 348 -84 349 -83
rect 349 -84 350 -83
rect 350 -84 351 -83
rect 351 -84 352 -83
rect 352 -84 353 -83
rect 353 -84 354 -83
rect 354 -84 355 -83
rect 355 -84 356 -83
rect 356 -84 357 -83
rect 357 -84 358 -83
rect 358 -84 359 -83
rect 359 -84 360 -83
rect 360 -84 361 -83
rect 361 -84 362 -83
rect 362 -84 363 -83
rect 363 -84 364 -83
rect 364 -84 365 -83
rect 365 -84 366 -83
rect 366 -84 367 -83
rect 367 -84 368 -83
rect 368 -84 369 -83
rect 369 -84 370 -83
rect 370 -84 371 -83
rect 371 -84 372 -83
rect 372 -84 373 -83
rect 373 -84 374 -83
rect 374 -84 375 -83
rect 375 -84 376 -83
rect 376 -84 377 -83
rect 377 -84 378 -83
rect 378 -84 379 -83
rect 379 -84 380 -83
rect 380 -84 381 -83
rect 381 -84 382 -83
rect 382 -84 383 -83
rect 383 -84 384 -83
rect 384 -84 385 -83
rect 385 -84 386 -83
rect 386 -84 387 -83
rect 387 -84 388 -83
rect 388 -84 389 -83
rect 389 -84 390 -83
rect 390 -84 391 -83
rect 391 -84 392 -83
rect 392 -84 393 -83
rect 393 -84 394 -83
rect 394 -84 395 -83
rect 395 -84 396 -83
rect 396 -84 397 -83
rect 397 -84 398 -83
rect 398 -84 399 -83
rect 399 -84 400 -83
rect 400 -84 401 -83
rect 401 -84 402 -83
rect 402 -84 403 -83
rect 403 -84 404 -83
rect 404 -84 405 -83
rect 405 -84 406 -83
rect 406 -84 407 -83
rect 407 -84 408 -83
rect 408 -84 409 -83
rect 409 -84 410 -83
rect 410 -84 411 -83
rect 411 -84 412 -83
rect 412 -84 413 -83
rect 413 -84 414 -83
rect 414 -84 415 -83
rect 415 -84 416 -83
rect 416 -84 417 -83
rect 417 -84 418 -83
rect 418 -84 419 -83
rect 419 -84 420 -83
rect 420 -84 421 -83
rect 421 -84 422 -83
rect 422 -84 423 -83
rect 423 -84 424 -83
rect 424 -84 425 -83
rect 425 -84 426 -83
rect 426 -84 427 -83
rect 427 -84 428 -83
rect 428 -84 429 -83
rect 429 -84 430 -83
rect 430 -84 431 -83
rect 431 -84 432 -83
rect 432 -84 433 -83
rect 433 -84 434 -83
rect 434 -84 435 -83
rect 435 -84 436 -83
rect 436 -84 437 -83
rect 437 -84 438 -83
rect 438 -84 439 -83
rect 439 -84 440 -83
rect 440 -84 441 -83
rect 441 -84 442 -83
rect 442 -84 443 -83
rect 443 -84 444 -83
rect 444 -84 445 -83
rect 445 -84 446 -83
rect 446 -84 447 -83
rect 447 -84 448 -83
rect 448 -84 449 -83
rect 449 -84 450 -83
rect 450 -84 451 -83
rect 451 -84 452 -83
rect 452 -84 453 -83
rect 453 -84 454 -83
rect 454 -84 455 -83
rect 455 -84 456 -83
rect 456 -84 457 -83
rect 457 -84 458 -83
rect 458 -84 459 -83
rect 459 -84 460 -83
rect 460 -84 461 -83
rect 461 -84 462 -83
rect 462 -84 463 -83
rect 463 -84 464 -83
rect 464 -84 465 -83
rect 465 -84 466 -83
rect 466 -84 467 -83
rect 467 -84 468 -83
rect 468 -84 469 -83
rect 469 -84 470 -83
rect 470 -84 471 -83
rect 471 -84 472 -83
rect 472 -84 473 -83
rect 473 -84 474 -83
rect 474 -84 475 -83
rect 475 -84 476 -83
rect 476 -84 477 -83
rect 477 -84 478 -83
rect 478 -84 479 -83
rect 479 -84 480 -83
rect 2 -85 3 -84
rect 3 -85 4 -84
rect 4 -85 5 -84
rect 5 -85 6 -84
rect 6 -85 7 -84
rect 7 -85 8 -84
rect 8 -85 9 -84
rect 9 -85 10 -84
rect 10 -85 11 -84
rect 11 -85 12 -84
rect 12 -85 13 -84
rect 13 -85 14 -84
rect 14 -85 15 -84
rect 15 -85 16 -84
rect 16 -85 17 -84
rect 17 -85 18 -84
rect 18 -85 19 -84
rect 19 -85 20 -84
rect 20 -85 21 -84
rect 21 -85 22 -84
rect 22 -85 23 -84
rect 23 -85 24 -84
rect 24 -85 25 -84
rect 25 -85 26 -84
rect 26 -85 27 -84
rect 27 -85 28 -84
rect 37 -85 38 -84
rect 38 -85 39 -84
rect 39 -85 40 -84
rect 40 -85 41 -84
rect 41 -85 42 -84
rect 42 -85 43 -84
rect 43 -85 44 -84
rect 44 -85 45 -84
rect 45 -85 46 -84
rect 46 -85 47 -84
rect 47 -85 48 -84
rect 48 -85 49 -84
rect 49 -85 50 -84
rect 50 -85 51 -84
rect 51 -85 52 -84
rect 52 -85 53 -84
rect 53 -85 54 -84
rect 54 -85 55 -84
rect 55 -85 56 -84
rect 56 -85 57 -84
rect 57 -85 58 -84
rect 58 -85 59 -84
rect 59 -85 60 -84
rect 69 -85 70 -84
rect 70 -85 71 -84
rect 71 -85 72 -84
rect 72 -85 73 -84
rect 73 -85 74 -84
rect 74 -85 75 -84
rect 75 -85 76 -84
rect 76 -85 77 -84
rect 77 -85 78 -84
rect 78 -85 79 -84
rect 79 -85 80 -84
rect 80 -85 81 -84
rect 81 -85 82 -84
rect 82 -85 83 -84
rect 83 -85 84 -84
rect 84 -85 85 -84
rect 85 -85 86 -84
rect 86 -85 87 -84
rect 87 -85 88 -84
rect 88 -85 89 -84
rect 89 -85 90 -84
rect 90 -85 91 -84
rect 91 -85 92 -84
rect 101 -85 102 -84
rect 102 -85 103 -84
rect 103 -85 104 -84
rect 104 -85 105 -84
rect 105 -85 106 -84
rect 106 -85 107 -84
rect 107 -85 108 -84
rect 108 -85 109 -84
rect 109 -85 110 -84
rect 110 -85 111 -84
rect 111 -85 112 -84
rect 112 -85 113 -84
rect 113 -85 114 -84
rect 114 -85 115 -84
rect 115 -85 116 -84
rect 116 -85 117 -84
rect 117 -85 118 -84
rect 118 -85 119 -84
rect 119 -85 120 -84
rect 120 -85 121 -84
rect 121 -85 122 -84
rect 122 -85 123 -84
rect 123 -85 124 -84
rect 133 -85 134 -84
rect 134 -85 135 -84
rect 135 -85 136 -84
rect 136 -85 137 -84
rect 137 -85 138 -84
rect 138 -85 139 -84
rect 139 -85 140 -84
rect 140 -85 141 -84
rect 141 -85 142 -84
rect 142 -85 143 -84
rect 143 -85 144 -84
rect 144 -85 145 -84
rect 145 -85 146 -84
rect 146 -85 147 -84
rect 147 -85 148 -84
rect 148 -85 149 -84
rect 149 -85 150 -84
rect 150 -85 151 -84
rect 151 -85 152 -84
rect 152 -85 153 -84
rect 153 -85 154 -84
rect 154 -85 155 -84
rect 155 -85 156 -84
rect 165 -85 166 -84
rect 166 -85 167 -84
rect 167 -85 168 -84
rect 168 -85 169 -84
rect 169 -85 170 -84
rect 170 -85 171 -84
rect 171 -85 172 -84
rect 172 -85 173 -84
rect 173 -85 174 -84
rect 174 -85 175 -84
rect 175 -85 176 -84
rect 176 -85 177 -84
rect 177 -85 178 -84
rect 178 -85 179 -84
rect 179 -85 180 -84
rect 180 -85 181 -84
rect 181 -85 182 -84
rect 182 -85 183 -84
rect 183 -85 184 -84
rect 184 -85 185 -84
rect 185 -85 186 -84
rect 186 -85 187 -84
rect 187 -85 188 -84
rect 188 -85 189 -84
rect 189 -85 190 -84
rect 190 -85 191 -84
rect 191 -85 192 -84
rect 192 -85 193 -84
rect 193 -85 194 -84
rect 194 -85 195 -84
rect 195 -85 196 -84
rect 196 -85 197 -84
rect 197 -85 198 -84
rect 198 -85 199 -84
rect 199 -85 200 -84
rect 200 -85 201 -84
rect 201 -85 202 -84
rect 202 -85 203 -84
rect 203 -85 204 -84
rect 204 -85 205 -84
rect 205 -85 206 -84
rect 206 -85 207 -84
rect 207 -85 208 -84
rect 208 -85 209 -84
rect 209 -85 210 -84
rect 210 -85 211 -84
rect 211 -85 212 -84
rect 212 -85 213 -84
rect 213 -85 214 -84
rect 214 -85 215 -84
rect 215 -85 216 -84
rect 216 -85 217 -84
rect 217 -85 218 -84
rect 218 -85 219 -84
rect 219 -85 220 -84
rect 220 -85 221 -84
rect 221 -85 222 -84
rect 222 -85 223 -84
rect 223 -85 224 -84
rect 224 -85 225 -84
rect 225 -85 226 -84
rect 226 -85 227 -84
rect 227 -85 228 -84
rect 228 -85 229 -84
rect 229 -85 230 -84
rect 230 -85 231 -84
rect 231 -85 232 -84
rect 232 -85 233 -84
rect 233 -85 234 -84
rect 234 -85 235 -84
rect 235 -85 236 -84
rect 236 -85 237 -84
rect 237 -85 238 -84
rect 238 -85 239 -84
rect 239 -85 240 -84
rect 240 -85 241 -84
rect 241 -85 242 -84
rect 242 -85 243 -84
rect 243 -85 244 -84
rect 244 -85 245 -84
rect 245 -85 246 -84
rect 246 -85 247 -84
rect 247 -85 248 -84
rect 248 -85 249 -84
rect 249 -85 250 -84
rect 250 -85 251 -84
rect 251 -85 252 -84
rect 252 -85 253 -84
rect 253 -85 254 -84
rect 254 -85 255 -84
rect 255 -85 256 -84
rect 256 -85 257 -84
rect 257 -85 258 -84
rect 258 -85 259 -84
rect 259 -85 260 -84
rect 260 -85 261 -84
rect 261 -85 262 -84
rect 262 -85 263 -84
rect 263 -85 264 -84
rect 264 -85 265 -84
rect 265 -85 266 -84
rect 266 -85 267 -84
rect 267 -85 268 -84
rect 268 -85 269 -84
rect 269 -85 270 -84
rect 270 -85 271 -84
rect 271 -85 272 -84
rect 272 -85 273 -84
rect 273 -85 274 -84
rect 274 -85 275 -84
rect 275 -85 276 -84
rect 276 -85 277 -84
rect 277 -85 278 -84
rect 278 -85 279 -84
rect 279 -85 280 -84
rect 280 -85 281 -84
rect 281 -85 282 -84
rect 282 -85 283 -84
rect 283 -85 284 -84
rect 284 -85 285 -84
rect 285 -85 286 -84
rect 286 -85 287 -84
rect 287 -85 288 -84
rect 288 -85 289 -84
rect 289 -85 290 -84
rect 290 -85 291 -84
rect 291 -85 292 -84
rect 292 -85 293 -84
rect 293 -85 294 -84
rect 294 -85 295 -84
rect 295 -85 296 -84
rect 296 -85 297 -84
rect 297 -85 298 -84
rect 298 -85 299 -84
rect 299 -85 300 -84
rect 300 -85 301 -84
rect 301 -85 302 -84
rect 302 -85 303 -84
rect 303 -85 304 -84
rect 304 -85 305 -84
rect 305 -85 306 -84
rect 306 -85 307 -84
rect 307 -85 308 -84
rect 308 -85 309 -84
rect 309 -85 310 -84
rect 310 -85 311 -84
rect 311 -85 312 -84
rect 312 -85 313 -84
rect 313 -85 314 -84
rect 314 -85 315 -84
rect 315 -85 316 -84
rect 316 -85 317 -84
rect 317 -85 318 -84
rect 318 -85 319 -84
rect 319 -85 320 -84
rect 320 -85 321 -84
rect 321 -85 322 -84
rect 322 -85 323 -84
rect 323 -85 324 -84
rect 324 -85 325 -84
rect 325 -85 326 -84
rect 326 -85 327 -84
rect 327 -85 328 -84
rect 328 -85 329 -84
rect 329 -85 330 -84
rect 330 -85 331 -84
rect 331 -85 332 -84
rect 332 -85 333 -84
rect 333 -85 334 -84
rect 334 -85 335 -84
rect 335 -85 336 -84
rect 336 -85 337 -84
rect 337 -85 338 -84
rect 338 -85 339 -84
rect 339 -85 340 -84
rect 340 -85 341 -84
rect 341 -85 342 -84
rect 342 -85 343 -84
rect 343 -85 344 -84
rect 344 -85 345 -84
rect 345 -85 346 -84
rect 346 -85 347 -84
rect 347 -85 348 -84
rect 348 -85 349 -84
rect 349 -85 350 -84
rect 350 -85 351 -84
rect 351 -85 352 -84
rect 352 -85 353 -84
rect 353 -85 354 -84
rect 354 -85 355 -84
rect 355 -85 356 -84
rect 356 -85 357 -84
rect 357 -85 358 -84
rect 358 -85 359 -84
rect 359 -85 360 -84
rect 360 -85 361 -84
rect 361 -85 362 -84
rect 362 -85 363 -84
rect 363 -85 364 -84
rect 364 -85 365 -84
rect 365 -85 366 -84
rect 366 -85 367 -84
rect 367 -85 368 -84
rect 368 -85 369 -84
rect 369 -85 370 -84
rect 370 -85 371 -84
rect 371 -85 372 -84
rect 372 -85 373 -84
rect 373 -85 374 -84
rect 374 -85 375 -84
rect 375 -85 376 -84
rect 376 -85 377 -84
rect 377 -85 378 -84
rect 378 -85 379 -84
rect 379 -85 380 -84
rect 380 -85 381 -84
rect 381 -85 382 -84
rect 382 -85 383 -84
rect 383 -85 384 -84
rect 384 -85 385 -84
rect 385 -85 386 -84
rect 386 -85 387 -84
rect 387 -85 388 -84
rect 388 -85 389 -84
rect 389 -85 390 -84
rect 390 -85 391 -84
rect 391 -85 392 -84
rect 392 -85 393 -84
rect 393 -85 394 -84
rect 394 -85 395 -84
rect 395 -85 396 -84
rect 396 -85 397 -84
rect 397 -85 398 -84
rect 398 -85 399 -84
rect 399 -85 400 -84
rect 400 -85 401 -84
rect 401 -85 402 -84
rect 402 -85 403 -84
rect 403 -85 404 -84
rect 404 -85 405 -84
rect 405 -85 406 -84
rect 406 -85 407 -84
rect 407 -85 408 -84
rect 408 -85 409 -84
rect 409 -85 410 -84
rect 410 -85 411 -84
rect 411 -85 412 -84
rect 412 -85 413 -84
rect 413 -85 414 -84
rect 414 -85 415 -84
rect 415 -85 416 -84
rect 416 -85 417 -84
rect 417 -85 418 -84
rect 418 -85 419 -84
rect 419 -85 420 -84
rect 420 -85 421 -84
rect 421 -85 422 -84
rect 422 -85 423 -84
rect 423 -85 424 -84
rect 424 -85 425 -84
rect 425 -85 426 -84
rect 426 -85 427 -84
rect 427 -85 428 -84
rect 428 -85 429 -84
rect 429 -85 430 -84
rect 430 -85 431 -84
rect 431 -85 432 -84
rect 432 -85 433 -84
rect 433 -85 434 -84
rect 434 -85 435 -84
rect 435 -85 436 -84
rect 436 -85 437 -84
rect 437 -85 438 -84
rect 438 -85 439 -84
rect 439 -85 440 -84
rect 440 -85 441 -84
rect 441 -85 442 -84
rect 442 -85 443 -84
rect 443 -85 444 -84
rect 444 -85 445 -84
rect 445 -85 446 -84
rect 446 -85 447 -84
rect 447 -85 448 -84
rect 448 -85 449 -84
rect 449 -85 450 -84
rect 450 -85 451 -84
rect 451 -85 452 -84
rect 452 -85 453 -84
rect 453 -85 454 -84
rect 454 -85 455 -84
rect 455 -85 456 -84
rect 456 -85 457 -84
rect 457 -85 458 -84
rect 458 -85 459 -84
rect 459 -85 460 -84
rect 460 -85 461 -84
rect 461 -85 462 -84
rect 462 -85 463 -84
rect 463 -85 464 -84
rect 464 -85 465 -84
rect 465 -85 466 -84
rect 466 -85 467 -84
rect 467 -85 468 -84
rect 468 -85 469 -84
rect 469 -85 470 -84
rect 470 -85 471 -84
rect 471 -85 472 -84
rect 472 -85 473 -84
rect 473 -85 474 -84
rect 474 -85 475 -84
rect 475 -85 476 -84
rect 476 -85 477 -84
rect 477 -85 478 -84
rect 478 -85 479 -84
rect 479 -85 480 -84
rect 2 -86 3 -85
rect 3 -86 4 -85
rect 4 -86 5 -85
rect 5 -86 6 -85
rect 6 -86 7 -85
rect 7 -86 8 -85
rect 8 -86 9 -85
rect 9 -86 10 -85
rect 10 -86 11 -85
rect 11 -86 12 -85
rect 12 -86 13 -85
rect 13 -86 14 -85
rect 14 -86 15 -85
rect 15 -86 16 -85
rect 16 -86 17 -85
rect 17 -86 18 -85
rect 18 -86 19 -85
rect 19 -86 20 -85
rect 20 -86 21 -85
rect 21 -86 22 -85
rect 22 -86 23 -85
rect 23 -86 24 -85
rect 24 -86 25 -85
rect 25 -86 26 -85
rect 26 -86 27 -85
rect 27 -86 28 -85
rect 32 -86 33 -85
rect 38 -86 39 -85
rect 39 -86 40 -85
rect 40 -86 41 -85
rect 41 -86 42 -85
rect 42 -86 43 -85
rect 43 -86 44 -85
rect 44 -86 45 -85
rect 45 -86 46 -85
rect 46 -86 47 -85
rect 47 -86 48 -85
rect 48 -86 49 -85
rect 49 -86 50 -85
rect 50 -86 51 -85
rect 51 -86 52 -85
rect 52 -86 53 -85
rect 53 -86 54 -85
rect 54 -86 55 -85
rect 55 -86 56 -85
rect 56 -86 57 -85
rect 57 -86 58 -85
rect 58 -86 59 -85
rect 59 -86 60 -85
rect 64 -86 65 -85
rect 69 -86 70 -85
rect 70 -86 71 -85
rect 71 -86 72 -85
rect 72 -86 73 -85
rect 73 -86 74 -85
rect 74 -86 75 -85
rect 75 -86 76 -85
rect 76 -86 77 -85
rect 77 -86 78 -85
rect 78 -86 79 -85
rect 79 -86 80 -85
rect 80 -86 81 -85
rect 81 -86 82 -85
rect 82 -86 83 -85
rect 83 -86 84 -85
rect 84 -86 85 -85
rect 85 -86 86 -85
rect 86 -86 87 -85
rect 87 -86 88 -85
rect 88 -86 89 -85
rect 89 -86 90 -85
rect 90 -86 91 -85
rect 91 -86 92 -85
rect 96 -86 97 -85
rect 102 -86 103 -85
rect 103 -86 104 -85
rect 104 -86 105 -85
rect 105 -86 106 -85
rect 106 -86 107 -85
rect 107 -86 108 -85
rect 108 -86 109 -85
rect 109 -86 110 -85
rect 110 -86 111 -85
rect 111 -86 112 -85
rect 112 -86 113 -85
rect 113 -86 114 -85
rect 114 -86 115 -85
rect 115 -86 116 -85
rect 116 -86 117 -85
rect 117 -86 118 -85
rect 118 -86 119 -85
rect 119 -86 120 -85
rect 120 -86 121 -85
rect 121 -86 122 -85
rect 122 -86 123 -85
rect 123 -86 124 -85
rect 128 -86 129 -85
rect 133 -86 134 -85
rect 134 -86 135 -85
rect 135 -86 136 -85
rect 136 -86 137 -85
rect 137 -86 138 -85
rect 138 -86 139 -85
rect 139 -86 140 -85
rect 140 -86 141 -85
rect 141 -86 142 -85
rect 142 -86 143 -85
rect 143 -86 144 -85
rect 144 -86 145 -85
rect 145 -86 146 -85
rect 146 -86 147 -85
rect 147 -86 148 -85
rect 148 -86 149 -85
rect 149 -86 150 -85
rect 150 -86 151 -85
rect 151 -86 152 -85
rect 152 -86 153 -85
rect 153 -86 154 -85
rect 154 -86 155 -85
rect 155 -86 156 -85
rect 160 -86 161 -85
rect 166 -86 167 -85
rect 167 -86 168 -85
rect 168 -86 169 -85
rect 169 -86 170 -85
rect 170 -86 171 -85
rect 171 -86 172 -85
rect 172 -86 173 -85
rect 173 -86 174 -85
rect 174 -86 175 -85
rect 175 -86 176 -85
rect 176 -86 177 -85
rect 177 -86 178 -85
rect 178 -86 179 -85
rect 179 -86 180 -85
rect 180 -86 181 -85
rect 181 -86 182 -85
rect 182 -86 183 -85
rect 183 -86 184 -85
rect 184 -86 185 -85
rect 185 -86 186 -85
rect 186 -86 187 -85
rect 187 -86 188 -85
rect 188 -86 189 -85
rect 189 -86 190 -85
rect 190 -86 191 -85
rect 191 -86 192 -85
rect 192 -86 193 -85
rect 193 -86 194 -85
rect 194 -86 195 -85
rect 195 -86 196 -85
rect 196 -86 197 -85
rect 197 -86 198 -85
rect 198 -86 199 -85
rect 199 -86 200 -85
rect 200 -86 201 -85
rect 201 -86 202 -85
rect 202 -86 203 -85
rect 203 -86 204 -85
rect 204 -86 205 -85
rect 205 -86 206 -85
rect 206 -86 207 -85
rect 207 -86 208 -85
rect 208 -86 209 -85
rect 209 -86 210 -85
rect 210 -86 211 -85
rect 211 -86 212 -85
rect 212 -86 213 -85
rect 213 -86 214 -85
rect 214 -86 215 -85
rect 215 -86 216 -85
rect 216 -86 217 -85
rect 217 -86 218 -85
rect 218 -86 219 -85
rect 219 -86 220 -85
rect 220 -86 221 -85
rect 221 -86 222 -85
rect 222 -86 223 -85
rect 223 -86 224 -85
rect 224 -86 225 -85
rect 225 -86 226 -85
rect 226 -86 227 -85
rect 227 -86 228 -85
rect 228 -86 229 -85
rect 229 -86 230 -85
rect 230 -86 231 -85
rect 231 -86 232 -85
rect 232 -86 233 -85
rect 233 -86 234 -85
rect 234 -86 235 -85
rect 235 -86 236 -85
rect 236 -86 237 -85
rect 237 -86 238 -85
rect 238 -86 239 -85
rect 239 -86 240 -85
rect 240 -86 241 -85
rect 241 -86 242 -85
rect 242 -86 243 -85
rect 243 -86 244 -85
rect 244 -86 245 -85
rect 245 -86 246 -85
rect 246 -86 247 -85
rect 247 -86 248 -85
rect 248 -86 249 -85
rect 249 -86 250 -85
rect 250 -86 251 -85
rect 251 -86 252 -85
rect 252 -86 253 -85
rect 253 -86 254 -85
rect 254 -86 255 -85
rect 255 -86 256 -85
rect 256 -86 257 -85
rect 257 -86 258 -85
rect 258 -86 259 -85
rect 259 -86 260 -85
rect 260 -86 261 -85
rect 261 -86 262 -85
rect 262 -86 263 -85
rect 263 -86 264 -85
rect 264 -86 265 -85
rect 265 -86 266 -85
rect 266 -86 267 -85
rect 267 -86 268 -85
rect 268 -86 269 -85
rect 269 -86 270 -85
rect 270 -86 271 -85
rect 271 -86 272 -85
rect 272 -86 273 -85
rect 273 -86 274 -85
rect 274 -86 275 -85
rect 275 -86 276 -85
rect 276 -86 277 -85
rect 277 -86 278 -85
rect 278 -86 279 -85
rect 279 -86 280 -85
rect 280 -86 281 -85
rect 281 -86 282 -85
rect 282 -86 283 -85
rect 283 -86 284 -85
rect 284 -86 285 -85
rect 285 -86 286 -85
rect 286 -86 287 -85
rect 287 -86 288 -85
rect 288 -86 289 -85
rect 289 -86 290 -85
rect 290 -86 291 -85
rect 291 -86 292 -85
rect 292 -86 293 -85
rect 293 -86 294 -85
rect 294 -86 295 -85
rect 295 -86 296 -85
rect 296 -86 297 -85
rect 297 -86 298 -85
rect 298 -86 299 -85
rect 299 -86 300 -85
rect 300 -86 301 -85
rect 301 -86 302 -85
rect 302 -86 303 -85
rect 303 -86 304 -85
rect 304 -86 305 -85
rect 305 -86 306 -85
rect 306 -86 307 -85
rect 307 -86 308 -85
rect 308 -86 309 -85
rect 309 -86 310 -85
rect 310 -86 311 -85
rect 311 -86 312 -85
rect 312 -86 313 -85
rect 313 -86 314 -85
rect 314 -86 315 -85
rect 315 -86 316 -85
rect 316 -86 317 -85
rect 317 -86 318 -85
rect 318 -86 319 -85
rect 319 -86 320 -85
rect 320 -86 321 -85
rect 321 -86 322 -85
rect 322 -86 323 -85
rect 323 -86 324 -85
rect 324 -86 325 -85
rect 325 -86 326 -85
rect 326 -86 327 -85
rect 327 -86 328 -85
rect 328 -86 329 -85
rect 329 -86 330 -85
rect 330 -86 331 -85
rect 331 -86 332 -85
rect 332 -86 333 -85
rect 333 -86 334 -85
rect 334 -86 335 -85
rect 335 -86 336 -85
rect 336 -86 337 -85
rect 337 -86 338 -85
rect 338 -86 339 -85
rect 339 -86 340 -85
rect 340 -86 341 -85
rect 341 -86 342 -85
rect 342 -86 343 -85
rect 343 -86 344 -85
rect 344 -86 345 -85
rect 345 -86 346 -85
rect 346 -86 347 -85
rect 347 -86 348 -85
rect 348 -86 349 -85
rect 349 -86 350 -85
rect 350 -86 351 -85
rect 351 -86 352 -85
rect 352 -86 353 -85
rect 353 -86 354 -85
rect 354 -86 355 -85
rect 355 -86 356 -85
rect 356 -86 357 -85
rect 357 -86 358 -85
rect 358 -86 359 -85
rect 359 -86 360 -85
rect 360 -86 361 -85
rect 361 -86 362 -85
rect 362 -86 363 -85
rect 363 -86 364 -85
rect 364 -86 365 -85
rect 365 -86 366 -85
rect 366 -86 367 -85
rect 367 -86 368 -85
rect 368 -86 369 -85
rect 369 -86 370 -85
rect 370 -86 371 -85
rect 371 -86 372 -85
rect 372 -86 373 -85
rect 373 -86 374 -85
rect 374 -86 375 -85
rect 375 -86 376 -85
rect 376 -86 377 -85
rect 377 -86 378 -85
rect 378 -86 379 -85
rect 379 -86 380 -85
rect 380 -86 381 -85
rect 381 -86 382 -85
rect 382 -86 383 -85
rect 383 -86 384 -85
rect 384 -86 385 -85
rect 385 -86 386 -85
rect 386 -86 387 -85
rect 387 -86 388 -85
rect 388 -86 389 -85
rect 389 -86 390 -85
rect 390 -86 391 -85
rect 391 -86 392 -85
rect 392 -86 393 -85
rect 393 -86 394 -85
rect 394 -86 395 -85
rect 395 -86 396 -85
rect 396 -86 397 -85
rect 397 -86 398 -85
rect 398 -86 399 -85
rect 399 -86 400 -85
rect 400 -86 401 -85
rect 401 -86 402 -85
rect 402 -86 403 -85
rect 403 -86 404 -85
rect 404 -86 405 -85
rect 405 -86 406 -85
rect 406 -86 407 -85
rect 407 -86 408 -85
rect 408 -86 409 -85
rect 409 -86 410 -85
rect 410 -86 411 -85
rect 411 -86 412 -85
rect 412 -86 413 -85
rect 413 -86 414 -85
rect 414 -86 415 -85
rect 415 -86 416 -85
rect 416 -86 417 -85
rect 417 -86 418 -85
rect 418 -86 419 -85
rect 419 -86 420 -85
rect 420 -86 421 -85
rect 421 -86 422 -85
rect 422 -86 423 -85
rect 423 -86 424 -85
rect 424 -86 425 -85
rect 425 -86 426 -85
rect 426 -86 427 -85
rect 427 -86 428 -85
rect 428 -86 429 -85
rect 429 -86 430 -85
rect 430 -86 431 -85
rect 431 -86 432 -85
rect 432 -86 433 -85
rect 433 -86 434 -85
rect 434 -86 435 -85
rect 435 -86 436 -85
rect 436 -86 437 -85
rect 437 -86 438 -85
rect 438 -86 439 -85
rect 439 -86 440 -85
rect 440 -86 441 -85
rect 441 -86 442 -85
rect 442 -86 443 -85
rect 443 -86 444 -85
rect 444 -86 445 -85
rect 445 -86 446 -85
rect 446 -86 447 -85
rect 447 -86 448 -85
rect 448 -86 449 -85
rect 449 -86 450 -85
rect 450 -86 451 -85
rect 451 -86 452 -85
rect 452 -86 453 -85
rect 453 -86 454 -85
rect 454 -86 455 -85
rect 455 -86 456 -85
rect 456 -86 457 -85
rect 457 -86 458 -85
rect 458 -86 459 -85
rect 459 -86 460 -85
rect 460 -86 461 -85
rect 461 -86 462 -85
rect 462 -86 463 -85
rect 463 -86 464 -85
rect 464 -86 465 -85
rect 465 -86 466 -85
rect 466 -86 467 -85
rect 467 -86 468 -85
rect 468 -86 469 -85
rect 469 -86 470 -85
rect 470 -86 471 -85
rect 471 -86 472 -85
rect 472 -86 473 -85
rect 473 -86 474 -85
rect 474 -86 475 -85
rect 475 -86 476 -85
rect 476 -86 477 -85
rect 477 -86 478 -85
rect 478 -86 479 -85
rect 479 -86 480 -85
rect 2 -87 3 -86
rect 3 -87 4 -86
rect 4 -87 5 -86
rect 5 -87 6 -86
rect 6 -87 7 -86
rect 7 -87 8 -86
rect 8 -87 9 -86
rect 9 -87 10 -86
rect 10 -87 11 -86
rect 11 -87 12 -86
rect 12 -87 13 -86
rect 13 -87 14 -86
rect 14 -87 15 -86
rect 15 -87 16 -86
rect 18 -87 19 -86
rect 19 -87 20 -86
rect 20 -87 21 -86
rect 21 -87 22 -86
rect 22 -87 23 -86
rect 23 -87 24 -86
rect 24 -87 25 -86
rect 25 -87 26 -86
rect 26 -87 27 -86
rect 27 -87 28 -86
rect 31 -87 32 -86
rect 32 -87 33 -86
rect 33 -87 34 -86
rect 34 -87 35 -86
rect 38 -87 39 -86
rect 39 -87 40 -86
rect 40 -87 41 -86
rect 41 -87 42 -86
rect 42 -87 43 -86
rect 43 -87 44 -86
rect 44 -87 45 -86
rect 45 -87 46 -86
rect 46 -87 47 -86
rect 47 -87 48 -86
rect 50 -87 51 -86
rect 51 -87 52 -86
rect 52 -87 53 -86
rect 53 -87 54 -86
rect 54 -87 55 -86
rect 55 -87 56 -86
rect 56 -87 57 -86
rect 57 -87 58 -86
rect 58 -87 59 -86
rect 59 -87 60 -86
rect 63 -87 64 -86
rect 64 -87 65 -86
rect 65 -87 66 -86
rect 69 -87 70 -86
rect 70 -87 71 -86
rect 71 -87 72 -86
rect 72 -87 73 -86
rect 73 -87 74 -86
rect 74 -87 75 -86
rect 75 -87 76 -86
rect 76 -87 77 -86
rect 77 -87 78 -86
rect 78 -87 79 -86
rect 79 -87 80 -86
rect 82 -87 83 -86
rect 83 -87 84 -86
rect 84 -87 85 -86
rect 85 -87 86 -86
rect 86 -87 87 -86
rect 87 -87 88 -86
rect 88 -87 89 -86
rect 89 -87 90 -86
rect 90 -87 91 -86
rect 91 -87 92 -86
rect 95 -87 96 -86
rect 96 -87 97 -86
rect 97 -87 98 -86
rect 98 -87 99 -86
rect 102 -87 103 -86
rect 103 -87 104 -86
rect 104 -87 105 -86
rect 105 -87 106 -86
rect 106 -87 107 -86
rect 107 -87 108 -86
rect 108 -87 109 -86
rect 109 -87 110 -86
rect 110 -87 111 -86
rect 111 -87 112 -86
rect 114 -87 115 -86
rect 115 -87 116 -86
rect 116 -87 117 -86
rect 117 -87 118 -86
rect 118 -87 119 -86
rect 119 -87 120 -86
rect 120 -87 121 -86
rect 121 -87 122 -86
rect 122 -87 123 -86
rect 123 -87 124 -86
rect 127 -87 128 -86
rect 128 -87 129 -86
rect 129 -87 130 -86
rect 133 -87 134 -86
rect 134 -87 135 -86
rect 135 -87 136 -86
rect 136 -87 137 -86
rect 137 -87 138 -86
rect 138 -87 139 -86
rect 139 -87 140 -86
rect 140 -87 141 -86
rect 141 -87 142 -86
rect 142 -87 143 -86
rect 143 -87 144 -86
rect 146 -87 147 -86
rect 147 -87 148 -86
rect 148 -87 149 -86
rect 149 -87 150 -86
rect 150 -87 151 -86
rect 151 -87 152 -86
rect 152 -87 153 -86
rect 153 -87 154 -86
rect 154 -87 155 -86
rect 155 -87 156 -86
rect 159 -87 160 -86
rect 160 -87 161 -86
rect 161 -87 162 -86
rect 162 -87 163 -86
rect 166 -87 167 -86
rect 167 -87 168 -86
rect 168 -87 169 -86
rect 169 -87 170 -86
rect 170 -87 171 -86
rect 171 -87 172 -86
rect 172 -87 173 -86
rect 173 -87 174 -86
rect 174 -87 175 -86
rect 175 -87 176 -86
rect 178 -87 179 -86
rect 179 -87 180 -86
rect 180 -87 181 -86
rect 181 -87 182 -86
rect 182 -87 183 -86
rect 183 -87 184 -86
rect 184 -87 185 -86
rect 185 -87 186 -86
rect 186 -87 187 -86
rect 187 -87 188 -86
rect 188 -87 189 -86
rect 189 -87 190 -86
rect 190 -87 191 -86
rect 191 -87 192 -86
rect 192 -87 193 -86
rect 193 -87 194 -86
rect 194 -87 195 -86
rect 195 -87 196 -86
rect 196 -87 197 -86
rect 197 -87 198 -86
rect 198 -87 199 -86
rect 199 -87 200 -86
rect 200 -87 201 -86
rect 201 -87 202 -86
rect 202 -87 203 -86
rect 203 -87 204 -86
rect 204 -87 205 -86
rect 205 -87 206 -86
rect 206 -87 207 -86
rect 207 -87 208 -86
rect 208 -87 209 -86
rect 209 -87 210 -86
rect 210 -87 211 -86
rect 211 -87 212 -86
rect 212 -87 213 -86
rect 213 -87 214 -86
rect 214 -87 215 -86
rect 215 -87 216 -86
rect 216 -87 217 -86
rect 217 -87 218 -86
rect 218 -87 219 -86
rect 219 -87 220 -86
rect 220 -87 221 -86
rect 221 -87 222 -86
rect 222 -87 223 -86
rect 223 -87 224 -86
rect 224 -87 225 -86
rect 225 -87 226 -86
rect 226 -87 227 -86
rect 227 -87 228 -86
rect 228 -87 229 -86
rect 229 -87 230 -86
rect 230 -87 231 -86
rect 231 -87 232 -86
rect 232 -87 233 -86
rect 233 -87 234 -86
rect 234 -87 235 -86
rect 235 -87 236 -86
rect 236 -87 237 -86
rect 237 -87 238 -86
rect 238 -87 239 -86
rect 239 -87 240 -86
rect 240 -87 241 -86
rect 241 -87 242 -86
rect 242 -87 243 -86
rect 243 -87 244 -86
rect 244 -87 245 -86
rect 245 -87 246 -86
rect 246 -87 247 -86
rect 247 -87 248 -86
rect 248 -87 249 -86
rect 249 -87 250 -86
rect 250 -87 251 -86
rect 251 -87 252 -86
rect 252 -87 253 -86
rect 253 -87 254 -86
rect 254 -87 255 -86
rect 255 -87 256 -86
rect 256 -87 257 -86
rect 257 -87 258 -86
rect 258 -87 259 -86
rect 259 -87 260 -86
rect 260 -87 261 -86
rect 261 -87 262 -86
rect 262 -87 263 -86
rect 263 -87 264 -86
rect 264 -87 265 -86
rect 265 -87 266 -86
rect 266 -87 267 -86
rect 267 -87 268 -86
rect 268 -87 269 -86
rect 269 -87 270 -86
rect 270 -87 271 -86
rect 271 -87 272 -86
rect 272 -87 273 -86
rect 273 -87 274 -86
rect 274 -87 275 -86
rect 275 -87 276 -86
rect 276 -87 277 -86
rect 277 -87 278 -86
rect 278 -87 279 -86
rect 279 -87 280 -86
rect 280 -87 281 -86
rect 281 -87 282 -86
rect 282 -87 283 -86
rect 283 -87 284 -86
rect 284 -87 285 -86
rect 285 -87 286 -86
rect 286 -87 287 -86
rect 287 -87 288 -86
rect 288 -87 289 -86
rect 289 -87 290 -86
rect 290 -87 291 -86
rect 291 -87 292 -86
rect 292 -87 293 -86
rect 293 -87 294 -86
rect 294 -87 295 -86
rect 295 -87 296 -86
rect 296 -87 297 -86
rect 297 -87 298 -86
rect 298 -87 299 -86
rect 299 -87 300 -86
rect 300 -87 301 -86
rect 301 -87 302 -86
rect 302 -87 303 -86
rect 303 -87 304 -86
rect 304 -87 305 -86
rect 305 -87 306 -86
rect 306 -87 307 -86
rect 307 -87 308 -86
rect 308 -87 309 -86
rect 309 -87 310 -86
rect 310 -87 311 -86
rect 311 -87 312 -86
rect 312 -87 313 -86
rect 313 -87 314 -86
rect 314 -87 315 -86
rect 315 -87 316 -86
rect 316 -87 317 -86
rect 317 -87 318 -86
rect 318 -87 319 -86
rect 319 -87 320 -86
rect 320 -87 321 -86
rect 321 -87 322 -86
rect 322 -87 323 -86
rect 323 -87 324 -86
rect 324 -87 325 -86
rect 325 -87 326 -86
rect 326 -87 327 -86
rect 327 -87 328 -86
rect 328 -87 329 -86
rect 329 -87 330 -86
rect 330 -87 331 -86
rect 331 -87 332 -86
rect 332 -87 333 -86
rect 333 -87 334 -86
rect 334 -87 335 -86
rect 335 -87 336 -86
rect 336 -87 337 -86
rect 337 -87 338 -86
rect 338 -87 339 -86
rect 339 -87 340 -86
rect 340 -87 341 -86
rect 341 -87 342 -86
rect 342 -87 343 -86
rect 343 -87 344 -86
rect 344 -87 345 -86
rect 345 -87 346 -86
rect 346 -87 347 -86
rect 347 -87 348 -86
rect 348 -87 349 -86
rect 349 -87 350 -86
rect 350 -87 351 -86
rect 351 -87 352 -86
rect 352 -87 353 -86
rect 353 -87 354 -86
rect 354 -87 355 -86
rect 355 -87 356 -86
rect 356 -87 357 -86
rect 357 -87 358 -86
rect 358 -87 359 -86
rect 359 -87 360 -86
rect 360 -87 361 -86
rect 361 -87 362 -86
rect 362 -87 363 -86
rect 363 -87 364 -86
rect 364 -87 365 -86
rect 365 -87 366 -86
rect 366 -87 367 -86
rect 367 -87 368 -86
rect 368 -87 369 -86
rect 369 -87 370 -86
rect 370 -87 371 -86
rect 371 -87 372 -86
rect 372 -87 373 -86
rect 373 -87 374 -86
rect 374 -87 375 -86
rect 375 -87 376 -86
rect 376 -87 377 -86
rect 377 -87 378 -86
rect 378 -87 379 -86
rect 379 -87 380 -86
rect 380 -87 381 -86
rect 381 -87 382 -86
rect 382 -87 383 -86
rect 383 -87 384 -86
rect 384 -87 385 -86
rect 385 -87 386 -86
rect 386 -87 387 -86
rect 387 -87 388 -86
rect 388 -87 389 -86
rect 389 -87 390 -86
rect 390 -87 391 -86
rect 391 -87 392 -86
rect 392 -87 393 -86
rect 393 -87 394 -86
rect 394 -87 395 -86
rect 395 -87 396 -86
rect 396 -87 397 -86
rect 397 -87 398 -86
rect 398 -87 399 -86
rect 399 -87 400 -86
rect 400 -87 401 -86
rect 401 -87 402 -86
rect 402 -87 403 -86
rect 403 -87 404 -86
rect 404 -87 405 -86
rect 405 -87 406 -86
rect 406 -87 407 -86
rect 407 -87 408 -86
rect 408 -87 409 -86
rect 409 -87 410 -86
rect 410 -87 411 -86
rect 411 -87 412 -86
rect 412 -87 413 -86
rect 413 -87 414 -86
rect 414 -87 415 -86
rect 415 -87 416 -86
rect 416 -87 417 -86
rect 417 -87 418 -86
rect 418 -87 419 -86
rect 419 -87 420 -86
rect 420 -87 421 -86
rect 421 -87 422 -86
rect 422 -87 423 -86
rect 423 -87 424 -86
rect 424 -87 425 -86
rect 425 -87 426 -86
rect 426 -87 427 -86
rect 427 -87 428 -86
rect 428 -87 429 -86
rect 429 -87 430 -86
rect 430 -87 431 -86
rect 431 -87 432 -86
rect 432 -87 433 -86
rect 433 -87 434 -86
rect 434 -87 435 -86
rect 435 -87 436 -86
rect 436 -87 437 -86
rect 437 -87 438 -86
rect 438 -87 439 -86
rect 439 -87 440 -86
rect 440 -87 441 -86
rect 441 -87 442 -86
rect 442 -87 443 -86
rect 443 -87 444 -86
rect 444 -87 445 -86
rect 445 -87 446 -86
rect 446 -87 447 -86
rect 447 -87 448 -86
rect 448 -87 449 -86
rect 449 -87 450 -86
rect 450 -87 451 -86
rect 451 -87 452 -86
rect 452 -87 453 -86
rect 453 -87 454 -86
rect 454 -87 455 -86
rect 455 -87 456 -86
rect 456 -87 457 -86
rect 457 -87 458 -86
rect 458 -87 459 -86
rect 459 -87 460 -86
rect 460 -87 461 -86
rect 461 -87 462 -86
rect 462 -87 463 -86
rect 463 -87 464 -86
rect 464 -87 465 -86
rect 465 -87 466 -86
rect 466 -87 467 -86
rect 467 -87 468 -86
rect 468 -87 469 -86
rect 469 -87 470 -86
rect 470 -87 471 -86
rect 471 -87 472 -86
rect 472 -87 473 -86
rect 473 -87 474 -86
rect 474 -87 475 -86
rect 475 -87 476 -86
rect 476 -87 477 -86
rect 477 -87 478 -86
rect 478 -87 479 -86
rect 479 -87 480 -86
rect 2 -88 3 -87
rect 3 -88 4 -87
rect 4 -88 5 -87
rect 5 -88 6 -87
rect 6 -88 7 -87
rect 7 -88 8 -87
rect 8 -88 9 -87
rect 9 -88 10 -87
rect 10 -88 11 -87
rect 11 -88 12 -87
rect 12 -88 13 -87
rect 13 -88 14 -87
rect 14 -88 15 -87
rect 18 -88 19 -87
rect 19 -88 20 -87
rect 20 -88 21 -87
rect 21 -88 22 -87
rect 22 -88 23 -87
rect 23 -88 24 -87
rect 24 -88 25 -87
rect 25 -88 26 -87
rect 26 -88 27 -87
rect 27 -88 28 -87
rect 30 -88 31 -87
rect 31 -88 32 -87
rect 32 -88 33 -87
rect 33 -88 34 -87
rect 34 -88 35 -87
rect 35 -88 36 -87
rect 38 -88 39 -87
rect 39 -88 40 -87
rect 40 -88 41 -87
rect 41 -88 42 -87
rect 42 -88 43 -87
rect 43 -88 44 -87
rect 44 -88 45 -87
rect 45 -88 46 -87
rect 46 -88 47 -87
rect 50 -88 51 -87
rect 51 -88 52 -87
rect 52 -88 53 -87
rect 53 -88 54 -87
rect 54 -88 55 -87
rect 55 -88 56 -87
rect 56 -88 57 -87
rect 57 -88 58 -87
rect 58 -88 59 -87
rect 59 -88 60 -87
rect 60 -88 61 -87
rect 61 -88 62 -87
rect 62 -88 63 -87
rect 63 -88 64 -87
rect 64 -88 65 -87
rect 65 -88 66 -87
rect 66 -88 67 -87
rect 67 -88 68 -87
rect 68 -88 69 -87
rect 69 -88 70 -87
rect 70 -88 71 -87
rect 71 -88 72 -87
rect 72 -88 73 -87
rect 73 -88 74 -87
rect 74 -88 75 -87
rect 75 -88 76 -87
rect 76 -88 77 -87
rect 77 -88 78 -87
rect 78 -88 79 -87
rect 82 -88 83 -87
rect 83 -88 84 -87
rect 84 -88 85 -87
rect 85 -88 86 -87
rect 86 -88 87 -87
rect 87 -88 88 -87
rect 88 -88 89 -87
rect 89 -88 90 -87
rect 90 -88 91 -87
rect 91 -88 92 -87
rect 94 -88 95 -87
rect 95 -88 96 -87
rect 96 -88 97 -87
rect 97 -88 98 -87
rect 98 -88 99 -87
rect 99 -88 100 -87
rect 102 -88 103 -87
rect 103 -88 104 -87
rect 104 -88 105 -87
rect 105 -88 106 -87
rect 106 -88 107 -87
rect 107 -88 108 -87
rect 108 -88 109 -87
rect 109 -88 110 -87
rect 110 -88 111 -87
rect 114 -88 115 -87
rect 115 -88 116 -87
rect 116 -88 117 -87
rect 117 -88 118 -87
rect 118 -88 119 -87
rect 119 -88 120 -87
rect 120 -88 121 -87
rect 121 -88 122 -87
rect 122 -88 123 -87
rect 123 -88 124 -87
rect 124 -88 125 -87
rect 125 -88 126 -87
rect 126 -88 127 -87
rect 127 -88 128 -87
rect 128 -88 129 -87
rect 129 -88 130 -87
rect 130 -88 131 -87
rect 131 -88 132 -87
rect 132 -88 133 -87
rect 133 -88 134 -87
rect 134 -88 135 -87
rect 135 -88 136 -87
rect 136 -88 137 -87
rect 137 -88 138 -87
rect 138 -88 139 -87
rect 139 -88 140 -87
rect 140 -88 141 -87
rect 141 -88 142 -87
rect 142 -88 143 -87
rect 146 -88 147 -87
rect 147 -88 148 -87
rect 148 -88 149 -87
rect 149 -88 150 -87
rect 150 -88 151 -87
rect 151 -88 152 -87
rect 152 -88 153 -87
rect 153 -88 154 -87
rect 154 -88 155 -87
rect 155 -88 156 -87
rect 158 -88 159 -87
rect 159 -88 160 -87
rect 160 -88 161 -87
rect 161 -88 162 -87
rect 162 -88 163 -87
rect 163 -88 164 -87
rect 166 -88 167 -87
rect 167 -88 168 -87
rect 168 -88 169 -87
rect 169 -88 170 -87
rect 170 -88 171 -87
rect 171 -88 172 -87
rect 172 -88 173 -87
rect 173 -88 174 -87
rect 174 -88 175 -87
rect 178 -88 179 -87
rect 179 -88 180 -87
rect 180 -88 181 -87
rect 181 -88 182 -87
rect 182 -88 183 -87
rect 183 -88 184 -87
rect 184 -88 185 -87
rect 185 -88 186 -87
rect 186 -88 187 -87
rect 187 -88 188 -87
rect 188 -88 189 -87
rect 189 -88 190 -87
rect 190 -88 191 -87
rect 191 -88 192 -87
rect 192 -88 193 -87
rect 193 -88 194 -87
rect 194 -88 195 -87
rect 195 -88 196 -87
rect 196 -88 197 -87
rect 197 -88 198 -87
rect 198 -88 199 -87
rect 199 -88 200 -87
rect 200 -88 201 -87
rect 201 -88 202 -87
rect 202 -88 203 -87
rect 203 -88 204 -87
rect 204 -88 205 -87
rect 205 -88 206 -87
rect 206 -88 207 -87
rect 207 -88 208 -87
rect 208 -88 209 -87
rect 209 -88 210 -87
rect 210 -88 211 -87
rect 211 -88 212 -87
rect 212 -88 213 -87
rect 213 -88 214 -87
rect 214 -88 215 -87
rect 215 -88 216 -87
rect 216 -88 217 -87
rect 217 -88 218 -87
rect 218 -88 219 -87
rect 219 -88 220 -87
rect 220 -88 221 -87
rect 221 -88 222 -87
rect 222 -88 223 -87
rect 223 -88 224 -87
rect 224 -88 225 -87
rect 225 -88 226 -87
rect 226 -88 227 -87
rect 227 -88 228 -87
rect 228 -88 229 -87
rect 229 -88 230 -87
rect 230 -88 231 -87
rect 231 -88 232 -87
rect 232 -88 233 -87
rect 233 -88 234 -87
rect 234 -88 235 -87
rect 235 -88 236 -87
rect 236 -88 237 -87
rect 237 -88 238 -87
rect 238 -88 239 -87
rect 239 -88 240 -87
rect 240 -88 241 -87
rect 241 -88 242 -87
rect 242 -88 243 -87
rect 243 -88 244 -87
rect 244 -88 245 -87
rect 245 -88 246 -87
rect 246 -88 247 -87
rect 247 -88 248 -87
rect 248 -88 249 -87
rect 249 -88 250 -87
rect 250 -88 251 -87
rect 251 -88 252 -87
rect 252 -88 253 -87
rect 253 -88 254 -87
rect 254 -88 255 -87
rect 255 -88 256 -87
rect 256 -88 257 -87
rect 257 -88 258 -87
rect 258 -88 259 -87
rect 259 -88 260 -87
rect 260 -88 261 -87
rect 261 -88 262 -87
rect 262 -88 263 -87
rect 263 -88 264 -87
rect 264 -88 265 -87
rect 265 -88 266 -87
rect 266 -88 267 -87
rect 267 -88 268 -87
rect 268 -88 269 -87
rect 269 -88 270 -87
rect 270 -88 271 -87
rect 271 -88 272 -87
rect 272 -88 273 -87
rect 273 -88 274 -87
rect 274 -88 275 -87
rect 275 -88 276 -87
rect 276 -88 277 -87
rect 277 -88 278 -87
rect 278 -88 279 -87
rect 279 -88 280 -87
rect 280 -88 281 -87
rect 281 -88 282 -87
rect 282 -88 283 -87
rect 283 -88 284 -87
rect 284 -88 285 -87
rect 285 -88 286 -87
rect 286 -88 287 -87
rect 287 -88 288 -87
rect 288 -88 289 -87
rect 289 -88 290 -87
rect 290 -88 291 -87
rect 291 -88 292 -87
rect 292 -88 293 -87
rect 293 -88 294 -87
rect 294 -88 295 -87
rect 295 -88 296 -87
rect 296 -88 297 -87
rect 297 -88 298 -87
rect 298 -88 299 -87
rect 299 -88 300 -87
rect 300 -88 301 -87
rect 301 -88 302 -87
rect 302 -88 303 -87
rect 303 -88 304 -87
rect 304 -88 305 -87
rect 305 -88 306 -87
rect 306 -88 307 -87
rect 307 -88 308 -87
rect 308 -88 309 -87
rect 309 -88 310 -87
rect 310 -88 311 -87
rect 311 -88 312 -87
rect 312 -88 313 -87
rect 313 -88 314 -87
rect 314 -88 315 -87
rect 315 -88 316 -87
rect 316 -88 317 -87
rect 317 -88 318 -87
rect 318 -88 319 -87
rect 319 -88 320 -87
rect 320 -88 321 -87
rect 321 -88 322 -87
rect 322 -88 323 -87
rect 323 -88 324 -87
rect 324 -88 325 -87
rect 325 -88 326 -87
rect 326 -88 327 -87
rect 327 -88 328 -87
rect 328 -88 329 -87
rect 329 -88 330 -87
rect 330 -88 331 -87
rect 331 -88 332 -87
rect 332 -88 333 -87
rect 333 -88 334 -87
rect 334 -88 335 -87
rect 335 -88 336 -87
rect 336 -88 337 -87
rect 337 -88 338 -87
rect 338 -88 339 -87
rect 339 -88 340 -87
rect 340 -88 341 -87
rect 341 -88 342 -87
rect 342 -88 343 -87
rect 343 -88 344 -87
rect 344 -88 345 -87
rect 345 -88 346 -87
rect 346 -88 347 -87
rect 347 -88 348 -87
rect 348 -88 349 -87
rect 349 -88 350 -87
rect 350 -88 351 -87
rect 351 -88 352 -87
rect 352 -88 353 -87
rect 353 -88 354 -87
rect 354 -88 355 -87
rect 355 -88 356 -87
rect 356 -88 357 -87
rect 357 -88 358 -87
rect 358 -88 359 -87
rect 359 -88 360 -87
rect 360 -88 361 -87
rect 361 -88 362 -87
rect 362 -88 363 -87
rect 363 -88 364 -87
rect 364 -88 365 -87
rect 365 -88 366 -87
rect 366 -88 367 -87
rect 367 -88 368 -87
rect 368 -88 369 -87
rect 369 -88 370 -87
rect 370 -88 371 -87
rect 371 -88 372 -87
rect 372 -88 373 -87
rect 373 -88 374 -87
rect 374 -88 375 -87
rect 375 -88 376 -87
rect 376 -88 377 -87
rect 377 -88 378 -87
rect 378 -88 379 -87
rect 379 -88 380 -87
rect 380 -88 381 -87
rect 381 -88 382 -87
rect 382 -88 383 -87
rect 383 -88 384 -87
rect 384 -88 385 -87
rect 385 -88 386 -87
rect 386 -88 387 -87
rect 387 -88 388 -87
rect 388 -88 389 -87
rect 389 -88 390 -87
rect 390 -88 391 -87
rect 391 -88 392 -87
rect 392 -88 393 -87
rect 393 -88 394 -87
rect 394 -88 395 -87
rect 395 -88 396 -87
rect 396 -88 397 -87
rect 397 -88 398 -87
rect 398 -88 399 -87
rect 399 -88 400 -87
rect 400 -88 401 -87
rect 401 -88 402 -87
rect 402 -88 403 -87
rect 403 -88 404 -87
rect 404 -88 405 -87
rect 405 -88 406 -87
rect 406 -88 407 -87
rect 407 -88 408 -87
rect 408 -88 409 -87
rect 409 -88 410 -87
rect 410 -88 411 -87
rect 411 -88 412 -87
rect 412 -88 413 -87
rect 413 -88 414 -87
rect 414 -88 415 -87
rect 415 -88 416 -87
rect 416 -88 417 -87
rect 417 -88 418 -87
rect 418 -88 419 -87
rect 419 -88 420 -87
rect 420 -88 421 -87
rect 421 -88 422 -87
rect 422 -88 423 -87
rect 423 -88 424 -87
rect 424 -88 425 -87
rect 425 -88 426 -87
rect 426 -88 427 -87
rect 427 -88 428 -87
rect 428 -88 429 -87
rect 429 -88 430 -87
rect 430 -88 431 -87
rect 431 -88 432 -87
rect 432 -88 433 -87
rect 433 -88 434 -87
rect 434 -88 435 -87
rect 435 -88 436 -87
rect 436 -88 437 -87
rect 437 -88 438 -87
rect 438 -88 439 -87
rect 439 -88 440 -87
rect 440 -88 441 -87
rect 441 -88 442 -87
rect 442 -88 443 -87
rect 443 -88 444 -87
rect 444 -88 445 -87
rect 445 -88 446 -87
rect 446 -88 447 -87
rect 447 -88 448 -87
rect 448 -88 449 -87
rect 449 -88 450 -87
rect 450 -88 451 -87
rect 451 -88 452 -87
rect 452 -88 453 -87
rect 453 -88 454 -87
rect 454 -88 455 -87
rect 455 -88 456 -87
rect 456 -88 457 -87
rect 457 -88 458 -87
rect 458 -88 459 -87
rect 459 -88 460 -87
rect 460 -88 461 -87
rect 461 -88 462 -87
rect 462 -88 463 -87
rect 463 -88 464 -87
rect 464 -88 465 -87
rect 465 -88 466 -87
rect 466 -88 467 -87
rect 467 -88 468 -87
rect 468 -88 469 -87
rect 469 -88 470 -87
rect 470 -88 471 -87
rect 471 -88 472 -87
rect 472 -88 473 -87
rect 473 -88 474 -87
rect 474 -88 475 -87
rect 475 -88 476 -87
rect 476 -88 477 -87
rect 477 -88 478 -87
rect 478 -88 479 -87
rect 479 -88 480 -87
rect 2 -89 3 -88
rect 3 -89 4 -88
rect 4 -89 5 -88
rect 5 -89 6 -88
rect 6 -89 7 -88
rect 7 -89 8 -88
rect 8 -89 9 -88
rect 9 -89 10 -88
rect 10 -89 11 -88
rect 11 -89 12 -88
rect 12 -89 13 -88
rect 13 -89 14 -88
rect 14 -89 15 -88
rect 18 -89 19 -88
rect 19 -89 20 -88
rect 20 -89 21 -88
rect 21 -89 22 -88
rect 22 -89 23 -88
rect 23 -89 24 -88
rect 24 -89 25 -88
rect 25 -89 26 -88
rect 26 -89 27 -88
rect 27 -89 28 -88
rect 28 -89 29 -88
rect 29 -89 30 -88
rect 30 -89 31 -88
rect 31 -89 32 -88
rect 32 -89 33 -88
rect 33 -89 34 -88
rect 34 -89 35 -88
rect 35 -89 36 -88
rect 36 -89 37 -88
rect 37 -89 38 -88
rect 38 -89 39 -88
rect 39 -89 40 -88
rect 40 -89 41 -88
rect 41 -89 42 -88
rect 42 -89 43 -88
rect 43 -89 44 -88
rect 44 -89 45 -88
rect 45 -89 46 -88
rect 46 -89 47 -88
rect 50 -89 51 -88
rect 51 -89 52 -88
rect 52 -89 53 -88
rect 53 -89 54 -88
rect 54 -89 55 -88
rect 55 -89 56 -88
rect 56 -89 57 -88
rect 57 -89 58 -88
rect 58 -89 59 -88
rect 59 -89 60 -88
rect 60 -89 61 -88
rect 61 -89 62 -88
rect 62 -89 63 -88
rect 63 -89 64 -88
rect 64 -89 65 -88
rect 65 -89 66 -88
rect 66 -89 67 -88
rect 67 -89 68 -88
rect 68 -89 69 -88
rect 69 -89 70 -88
rect 70 -89 71 -88
rect 71 -89 72 -88
rect 72 -89 73 -88
rect 73 -89 74 -88
rect 74 -89 75 -88
rect 75 -89 76 -88
rect 76 -89 77 -88
rect 77 -89 78 -88
rect 78 -89 79 -88
rect 82 -89 83 -88
rect 83 -89 84 -88
rect 84 -89 85 -88
rect 85 -89 86 -88
rect 86 -89 87 -88
rect 87 -89 88 -88
rect 88 -89 89 -88
rect 89 -89 90 -88
rect 90 -89 91 -88
rect 91 -89 92 -88
rect 92 -89 93 -88
rect 93 -89 94 -88
rect 94 -89 95 -88
rect 95 -89 96 -88
rect 96 -89 97 -88
rect 97 -89 98 -88
rect 98 -89 99 -88
rect 99 -89 100 -88
rect 100 -89 101 -88
rect 101 -89 102 -88
rect 102 -89 103 -88
rect 103 -89 104 -88
rect 104 -89 105 -88
rect 105 -89 106 -88
rect 106 -89 107 -88
rect 107 -89 108 -88
rect 108 -89 109 -88
rect 109 -89 110 -88
rect 110 -89 111 -88
rect 114 -89 115 -88
rect 115 -89 116 -88
rect 116 -89 117 -88
rect 117 -89 118 -88
rect 118 -89 119 -88
rect 119 -89 120 -88
rect 120 -89 121 -88
rect 121 -89 122 -88
rect 122 -89 123 -88
rect 123 -89 124 -88
rect 124 -89 125 -88
rect 125 -89 126 -88
rect 126 -89 127 -88
rect 127 -89 128 -88
rect 128 -89 129 -88
rect 129 -89 130 -88
rect 130 -89 131 -88
rect 131 -89 132 -88
rect 132 -89 133 -88
rect 133 -89 134 -88
rect 134 -89 135 -88
rect 135 -89 136 -88
rect 136 -89 137 -88
rect 137 -89 138 -88
rect 138 -89 139 -88
rect 139 -89 140 -88
rect 140 -89 141 -88
rect 141 -89 142 -88
rect 142 -89 143 -88
rect 146 -89 147 -88
rect 147 -89 148 -88
rect 148 -89 149 -88
rect 149 -89 150 -88
rect 150 -89 151 -88
rect 151 -89 152 -88
rect 152 -89 153 -88
rect 153 -89 154 -88
rect 154 -89 155 -88
rect 155 -89 156 -88
rect 156 -89 157 -88
rect 157 -89 158 -88
rect 158 -89 159 -88
rect 159 -89 160 -88
rect 160 -89 161 -88
rect 161 -89 162 -88
rect 162 -89 163 -88
rect 163 -89 164 -88
rect 164 -89 165 -88
rect 165 -89 166 -88
rect 166 -89 167 -88
rect 167 -89 168 -88
rect 168 -89 169 -88
rect 169 -89 170 -88
rect 170 -89 171 -88
rect 171 -89 172 -88
rect 172 -89 173 -88
rect 173 -89 174 -88
rect 174 -89 175 -88
rect 178 -89 179 -88
rect 179 -89 180 -88
rect 180 -89 181 -88
rect 181 -89 182 -88
rect 182 -89 183 -88
rect 183 -89 184 -88
rect 184 -89 185 -88
rect 185 -89 186 -88
rect 186 -89 187 -88
rect 187 -89 188 -88
rect 188 -89 189 -88
rect 189 -89 190 -88
rect 190 -89 191 -88
rect 191 -89 192 -88
rect 192 -89 193 -88
rect 193 -89 194 -88
rect 194 -89 195 -88
rect 195 -89 196 -88
rect 196 -89 197 -88
rect 197 -89 198 -88
rect 198 -89 199 -88
rect 199 -89 200 -88
rect 200 -89 201 -88
rect 201 -89 202 -88
rect 202 -89 203 -88
rect 203 -89 204 -88
rect 204 -89 205 -88
rect 205 -89 206 -88
rect 206 -89 207 -88
rect 207 -89 208 -88
rect 208 -89 209 -88
rect 209 -89 210 -88
rect 210 -89 211 -88
rect 211 -89 212 -88
rect 212 -89 213 -88
rect 213 -89 214 -88
rect 214 -89 215 -88
rect 215 -89 216 -88
rect 216 -89 217 -88
rect 217 -89 218 -88
rect 218 -89 219 -88
rect 219 -89 220 -88
rect 220 -89 221 -88
rect 221 -89 222 -88
rect 222 -89 223 -88
rect 223 -89 224 -88
rect 224 -89 225 -88
rect 225 -89 226 -88
rect 226 -89 227 -88
rect 227 -89 228 -88
rect 228 -89 229 -88
rect 229 -89 230 -88
rect 230 -89 231 -88
rect 231 -89 232 -88
rect 232 -89 233 -88
rect 233 -89 234 -88
rect 234 -89 235 -88
rect 235 -89 236 -88
rect 236 -89 237 -88
rect 237 -89 238 -88
rect 238 -89 239 -88
rect 239 -89 240 -88
rect 240 -89 241 -88
rect 241 -89 242 -88
rect 242 -89 243 -88
rect 243 -89 244 -88
rect 244 -89 245 -88
rect 245 -89 246 -88
rect 246 -89 247 -88
rect 247 -89 248 -88
rect 248 -89 249 -88
rect 249 -89 250 -88
rect 250 -89 251 -88
rect 251 -89 252 -88
rect 252 -89 253 -88
rect 253 -89 254 -88
rect 254 -89 255 -88
rect 255 -89 256 -88
rect 256 -89 257 -88
rect 257 -89 258 -88
rect 258 -89 259 -88
rect 259 -89 260 -88
rect 260 -89 261 -88
rect 261 -89 262 -88
rect 262 -89 263 -88
rect 263 -89 264 -88
rect 264 -89 265 -88
rect 265 -89 266 -88
rect 266 -89 267 -88
rect 267 -89 268 -88
rect 268 -89 269 -88
rect 269 -89 270 -88
rect 270 -89 271 -88
rect 271 -89 272 -88
rect 272 -89 273 -88
rect 273 -89 274 -88
rect 274 -89 275 -88
rect 275 -89 276 -88
rect 276 -89 277 -88
rect 277 -89 278 -88
rect 278 -89 279 -88
rect 279 -89 280 -88
rect 280 -89 281 -88
rect 281 -89 282 -88
rect 282 -89 283 -88
rect 283 -89 284 -88
rect 284 -89 285 -88
rect 285 -89 286 -88
rect 286 -89 287 -88
rect 287 -89 288 -88
rect 288 -89 289 -88
rect 289 -89 290 -88
rect 290 -89 291 -88
rect 291 -89 292 -88
rect 292 -89 293 -88
rect 293 -89 294 -88
rect 294 -89 295 -88
rect 295 -89 296 -88
rect 296 -89 297 -88
rect 297 -89 298 -88
rect 298 -89 299 -88
rect 299 -89 300 -88
rect 300 -89 301 -88
rect 301 -89 302 -88
rect 302 -89 303 -88
rect 303 -89 304 -88
rect 304 -89 305 -88
rect 305 -89 306 -88
rect 306 -89 307 -88
rect 307 -89 308 -88
rect 308 -89 309 -88
rect 309 -89 310 -88
rect 310 -89 311 -88
rect 311 -89 312 -88
rect 312 -89 313 -88
rect 313 -89 314 -88
rect 314 -89 315 -88
rect 315 -89 316 -88
rect 316 -89 317 -88
rect 317 -89 318 -88
rect 318 -89 319 -88
rect 319 -89 320 -88
rect 320 -89 321 -88
rect 321 -89 322 -88
rect 322 -89 323 -88
rect 323 -89 324 -88
rect 324 -89 325 -88
rect 325 -89 326 -88
rect 326 -89 327 -88
rect 327 -89 328 -88
rect 328 -89 329 -88
rect 329 -89 330 -88
rect 330 -89 331 -88
rect 331 -89 332 -88
rect 332 -89 333 -88
rect 333 -89 334 -88
rect 334 -89 335 -88
rect 335 -89 336 -88
rect 336 -89 337 -88
rect 337 -89 338 -88
rect 338 -89 339 -88
rect 339 -89 340 -88
rect 340 -89 341 -88
rect 341 -89 342 -88
rect 342 -89 343 -88
rect 343 -89 344 -88
rect 344 -89 345 -88
rect 345 -89 346 -88
rect 346 -89 347 -88
rect 347 -89 348 -88
rect 348 -89 349 -88
rect 349 -89 350 -88
rect 350 -89 351 -88
rect 351 -89 352 -88
rect 352 -89 353 -88
rect 353 -89 354 -88
rect 354 -89 355 -88
rect 355 -89 356 -88
rect 356 -89 357 -88
rect 357 -89 358 -88
rect 358 -89 359 -88
rect 359 -89 360 -88
rect 360 -89 361 -88
rect 361 -89 362 -88
rect 362 -89 363 -88
rect 363 -89 364 -88
rect 364 -89 365 -88
rect 365 -89 366 -88
rect 366 -89 367 -88
rect 367 -89 368 -88
rect 368 -89 369 -88
rect 369 -89 370 -88
rect 370 -89 371 -88
rect 371 -89 372 -88
rect 372 -89 373 -88
rect 373 -89 374 -88
rect 374 -89 375 -88
rect 375 -89 376 -88
rect 376 -89 377 -88
rect 377 -89 378 -88
rect 378 -89 379 -88
rect 379 -89 380 -88
rect 380 -89 381 -88
rect 381 -89 382 -88
rect 382 -89 383 -88
rect 383 -89 384 -88
rect 384 -89 385 -88
rect 385 -89 386 -88
rect 386 -89 387 -88
rect 387 -89 388 -88
rect 388 -89 389 -88
rect 389 -89 390 -88
rect 390 -89 391 -88
rect 391 -89 392 -88
rect 392 -89 393 -88
rect 393 -89 394 -88
rect 394 -89 395 -88
rect 395 -89 396 -88
rect 396 -89 397 -88
rect 397 -89 398 -88
rect 398 -89 399 -88
rect 399 -89 400 -88
rect 400 -89 401 -88
rect 401 -89 402 -88
rect 402 -89 403 -88
rect 403 -89 404 -88
rect 404 -89 405 -88
rect 405 -89 406 -88
rect 406 -89 407 -88
rect 407 -89 408 -88
rect 408 -89 409 -88
rect 409 -89 410 -88
rect 410 -89 411 -88
rect 411 -89 412 -88
rect 412 -89 413 -88
rect 413 -89 414 -88
rect 414 -89 415 -88
rect 415 -89 416 -88
rect 416 -89 417 -88
rect 417 -89 418 -88
rect 418 -89 419 -88
rect 419 -89 420 -88
rect 420 -89 421 -88
rect 421 -89 422 -88
rect 422 -89 423 -88
rect 423 -89 424 -88
rect 424 -89 425 -88
rect 425 -89 426 -88
rect 426 -89 427 -88
rect 427 -89 428 -88
rect 428 -89 429 -88
rect 429 -89 430 -88
rect 430 -89 431 -88
rect 431 -89 432 -88
rect 432 -89 433 -88
rect 433 -89 434 -88
rect 434 -89 435 -88
rect 435 -89 436 -88
rect 436 -89 437 -88
rect 437 -89 438 -88
rect 438 -89 439 -88
rect 439 -89 440 -88
rect 440 -89 441 -88
rect 441 -89 442 -88
rect 442 -89 443 -88
rect 443 -89 444 -88
rect 444 -89 445 -88
rect 445 -89 446 -88
rect 446 -89 447 -88
rect 447 -89 448 -88
rect 448 -89 449 -88
rect 449 -89 450 -88
rect 450 -89 451 -88
rect 451 -89 452 -88
rect 452 -89 453 -88
rect 453 -89 454 -88
rect 454 -89 455 -88
rect 455 -89 456 -88
rect 456 -89 457 -88
rect 457 -89 458 -88
rect 458 -89 459 -88
rect 459 -89 460 -88
rect 460 -89 461 -88
rect 461 -89 462 -88
rect 462 -89 463 -88
rect 463 -89 464 -88
rect 464 -89 465 -88
rect 465 -89 466 -88
rect 466 -89 467 -88
rect 467 -89 468 -88
rect 468 -89 469 -88
rect 469 -89 470 -88
rect 470 -89 471 -88
rect 471 -89 472 -88
rect 472 -89 473 -88
rect 473 -89 474 -88
rect 474 -89 475 -88
rect 475 -89 476 -88
rect 476 -89 477 -88
rect 477 -89 478 -88
rect 478 -89 479 -88
rect 479 -89 480 -88
rect 2 -90 3 -89
rect 3 -90 4 -89
rect 4 -90 5 -89
rect 5 -90 6 -89
rect 6 -90 7 -89
rect 7 -90 8 -89
rect 8 -90 9 -89
rect 9 -90 10 -89
rect 10 -90 11 -89
rect 11 -90 12 -89
rect 12 -90 13 -89
rect 13 -90 14 -89
rect 14 -90 15 -89
rect 19 -90 20 -89
rect 20 -90 21 -89
rect 21 -90 22 -89
rect 22 -90 23 -89
rect 23 -90 24 -89
rect 24 -90 25 -89
rect 25 -90 26 -89
rect 26 -90 27 -89
rect 27 -90 28 -89
rect 28 -90 29 -89
rect 29 -90 30 -89
rect 30 -90 31 -89
rect 31 -90 32 -89
rect 32 -90 33 -89
rect 33 -90 34 -89
rect 34 -90 35 -89
rect 35 -90 36 -89
rect 36 -90 37 -89
rect 37 -90 38 -89
rect 38 -90 39 -89
rect 39 -90 40 -89
rect 40 -90 41 -89
rect 41 -90 42 -89
rect 42 -90 43 -89
rect 43 -90 44 -89
rect 44 -90 45 -89
rect 45 -90 46 -89
rect 46 -90 47 -89
rect 51 -90 52 -89
rect 52 -90 53 -89
rect 53 -90 54 -89
rect 54 -90 55 -89
rect 55 -90 56 -89
rect 56 -90 57 -89
rect 57 -90 58 -89
rect 58 -90 59 -89
rect 59 -90 60 -89
rect 60 -90 61 -89
rect 61 -90 62 -89
rect 62 -90 63 -89
rect 63 -90 64 -89
rect 64 -90 65 -89
rect 65 -90 66 -89
rect 66 -90 67 -89
rect 67 -90 68 -89
rect 68 -90 69 -89
rect 69 -90 70 -89
rect 70 -90 71 -89
rect 71 -90 72 -89
rect 72 -90 73 -89
rect 73 -90 74 -89
rect 74 -90 75 -89
rect 75 -90 76 -89
rect 76 -90 77 -89
rect 77 -90 78 -89
rect 78 -90 79 -89
rect 83 -90 84 -89
rect 84 -90 85 -89
rect 85 -90 86 -89
rect 86 -90 87 -89
rect 87 -90 88 -89
rect 88 -90 89 -89
rect 89 -90 90 -89
rect 90 -90 91 -89
rect 91 -90 92 -89
rect 92 -90 93 -89
rect 93 -90 94 -89
rect 94 -90 95 -89
rect 95 -90 96 -89
rect 96 -90 97 -89
rect 97 -90 98 -89
rect 98 -90 99 -89
rect 99 -90 100 -89
rect 100 -90 101 -89
rect 101 -90 102 -89
rect 102 -90 103 -89
rect 103 -90 104 -89
rect 104 -90 105 -89
rect 105 -90 106 -89
rect 106 -90 107 -89
rect 107 -90 108 -89
rect 108 -90 109 -89
rect 109 -90 110 -89
rect 110 -90 111 -89
rect 115 -90 116 -89
rect 116 -90 117 -89
rect 117 -90 118 -89
rect 118 -90 119 -89
rect 119 -90 120 -89
rect 120 -90 121 -89
rect 121 -90 122 -89
rect 122 -90 123 -89
rect 123 -90 124 -89
rect 124 -90 125 -89
rect 125 -90 126 -89
rect 126 -90 127 -89
rect 127 -90 128 -89
rect 128 -90 129 -89
rect 129 -90 130 -89
rect 130 -90 131 -89
rect 131 -90 132 -89
rect 132 -90 133 -89
rect 133 -90 134 -89
rect 134 -90 135 -89
rect 135 -90 136 -89
rect 136 -90 137 -89
rect 137 -90 138 -89
rect 138 -90 139 -89
rect 139 -90 140 -89
rect 140 -90 141 -89
rect 141 -90 142 -89
rect 142 -90 143 -89
rect 147 -90 148 -89
rect 148 -90 149 -89
rect 149 -90 150 -89
rect 150 -90 151 -89
rect 151 -90 152 -89
rect 152 -90 153 -89
rect 153 -90 154 -89
rect 154 -90 155 -89
rect 155 -90 156 -89
rect 156 -90 157 -89
rect 157 -90 158 -89
rect 158 -90 159 -89
rect 159 -90 160 -89
rect 160 -90 161 -89
rect 161 -90 162 -89
rect 162 -90 163 -89
rect 163 -90 164 -89
rect 164 -90 165 -89
rect 165 -90 166 -89
rect 166 -90 167 -89
rect 167 -90 168 -89
rect 168 -90 169 -89
rect 169 -90 170 -89
rect 170 -90 171 -89
rect 171 -90 172 -89
rect 172 -90 173 -89
rect 173 -90 174 -89
rect 174 -90 175 -89
rect 179 -90 180 -89
rect 180 -90 181 -89
rect 181 -90 182 -89
rect 182 -90 183 -89
rect 183 -90 184 -89
rect 184 -90 185 -89
rect 185 -90 186 -89
rect 186 -90 187 -89
rect 187 -90 188 -89
rect 188 -90 189 -89
rect 189 -90 190 -89
rect 190 -90 191 -89
rect 191 -90 192 -89
rect 192 -90 193 -89
rect 193 -90 194 -89
rect 194 -90 195 -89
rect 195 -90 196 -89
rect 196 -90 197 -89
rect 197 -90 198 -89
rect 198 -90 199 -89
rect 199 -90 200 -89
rect 200 -90 201 -89
rect 201 -90 202 -89
rect 202 -90 203 -89
rect 203 -90 204 -89
rect 204 -90 205 -89
rect 205 -90 206 -89
rect 206 -90 207 -89
rect 207 -90 208 -89
rect 208 -90 209 -89
rect 209 -90 210 -89
rect 210 -90 211 -89
rect 211 -90 212 -89
rect 212 -90 213 -89
rect 213 -90 214 -89
rect 214 -90 215 -89
rect 215 -90 216 -89
rect 216 -90 217 -89
rect 217 -90 218 -89
rect 218 -90 219 -89
rect 219 -90 220 -89
rect 220 -90 221 -89
rect 221 -90 222 -89
rect 222 -90 223 -89
rect 223 -90 224 -89
rect 224 -90 225 -89
rect 225 -90 226 -89
rect 226 -90 227 -89
rect 227 -90 228 -89
rect 228 -90 229 -89
rect 229 -90 230 -89
rect 230 -90 231 -89
rect 231 -90 232 -89
rect 232 -90 233 -89
rect 233 -90 234 -89
rect 234 -90 235 -89
rect 235 -90 236 -89
rect 236 -90 237 -89
rect 237 -90 238 -89
rect 238 -90 239 -89
rect 239 -90 240 -89
rect 240 -90 241 -89
rect 241 -90 242 -89
rect 242 -90 243 -89
rect 243 -90 244 -89
rect 244 -90 245 -89
rect 245 -90 246 -89
rect 246 -90 247 -89
rect 247 -90 248 -89
rect 248 -90 249 -89
rect 249 -90 250 -89
rect 250 -90 251 -89
rect 251 -90 252 -89
rect 252 -90 253 -89
rect 253 -90 254 -89
rect 254 -90 255 -89
rect 255 -90 256 -89
rect 256 -90 257 -89
rect 257 -90 258 -89
rect 258 -90 259 -89
rect 259 -90 260 -89
rect 260 -90 261 -89
rect 261 -90 262 -89
rect 262 -90 263 -89
rect 263 -90 264 -89
rect 264 -90 265 -89
rect 265 -90 266 -89
rect 266 -90 267 -89
rect 267 -90 268 -89
rect 268 -90 269 -89
rect 269 -90 270 -89
rect 270 -90 271 -89
rect 271 -90 272 -89
rect 272 -90 273 -89
rect 273 -90 274 -89
rect 274 -90 275 -89
rect 275 -90 276 -89
rect 276 -90 277 -89
rect 277 -90 278 -89
rect 278 -90 279 -89
rect 279 -90 280 -89
rect 280 -90 281 -89
rect 281 -90 282 -89
rect 282 -90 283 -89
rect 283 -90 284 -89
rect 284 -90 285 -89
rect 285 -90 286 -89
rect 286 -90 287 -89
rect 287 -90 288 -89
rect 288 -90 289 -89
rect 289 -90 290 -89
rect 290 -90 291 -89
rect 291 -90 292 -89
rect 292 -90 293 -89
rect 293 -90 294 -89
rect 294 -90 295 -89
rect 295 -90 296 -89
rect 296 -90 297 -89
rect 297 -90 298 -89
rect 298 -90 299 -89
rect 299 -90 300 -89
rect 300 -90 301 -89
rect 301 -90 302 -89
rect 302 -90 303 -89
rect 303 -90 304 -89
rect 304 -90 305 -89
rect 305 -90 306 -89
rect 306 -90 307 -89
rect 307 -90 308 -89
rect 308 -90 309 -89
rect 309 -90 310 -89
rect 310 -90 311 -89
rect 311 -90 312 -89
rect 312 -90 313 -89
rect 313 -90 314 -89
rect 314 -90 315 -89
rect 315 -90 316 -89
rect 316 -90 317 -89
rect 317 -90 318 -89
rect 318 -90 319 -89
rect 319 -90 320 -89
rect 320 -90 321 -89
rect 321 -90 322 -89
rect 322 -90 323 -89
rect 323 -90 324 -89
rect 324 -90 325 -89
rect 325 -90 326 -89
rect 326 -90 327 -89
rect 327 -90 328 -89
rect 328 -90 329 -89
rect 329 -90 330 -89
rect 330 -90 331 -89
rect 331 -90 332 -89
rect 332 -90 333 -89
rect 333 -90 334 -89
rect 334 -90 335 -89
rect 335 -90 336 -89
rect 336 -90 337 -89
rect 337 -90 338 -89
rect 338 -90 339 -89
rect 339 -90 340 -89
rect 340 -90 341 -89
rect 341 -90 342 -89
rect 342 -90 343 -89
rect 343 -90 344 -89
rect 344 -90 345 -89
rect 345 -90 346 -89
rect 346 -90 347 -89
rect 347 -90 348 -89
rect 348 -90 349 -89
rect 349 -90 350 -89
rect 350 -90 351 -89
rect 351 -90 352 -89
rect 352 -90 353 -89
rect 353 -90 354 -89
rect 354 -90 355 -89
rect 355 -90 356 -89
rect 356 -90 357 -89
rect 357 -90 358 -89
rect 358 -90 359 -89
rect 359 -90 360 -89
rect 360 -90 361 -89
rect 361 -90 362 -89
rect 362 -90 363 -89
rect 363 -90 364 -89
rect 364 -90 365 -89
rect 365 -90 366 -89
rect 366 -90 367 -89
rect 367 -90 368 -89
rect 368 -90 369 -89
rect 369 -90 370 -89
rect 370 -90 371 -89
rect 371 -90 372 -89
rect 372 -90 373 -89
rect 373 -90 374 -89
rect 374 -90 375 -89
rect 375 -90 376 -89
rect 376 -90 377 -89
rect 377 -90 378 -89
rect 378 -90 379 -89
rect 379 -90 380 -89
rect 380 -90 381 -89
rect 381 -90 382 -89
rect 382 -90 383 -89
rect 383 -90 384 -89
rect 384 -90 385 -89
rect 385 -90 386 -89
rect 386 -90 387 -89
rect 387 -90 388 -89
rect 388 -90 389 -89
rect 389 -90 390 -89
rect 390 -90 391 -89
rect 391 -90 392 -89
rect 392 -90 393 -89
rect 393 -90 394 -89
rect 394 -90 395 -89
rect 395 -90 396 -89
rect 396 -90 397 -89
rect 397 -90 398 -89
rect 398 -90 399 -89
rect 399 -90 400 -89
rect 400 -90 401 -89
rect 401 -90 402 -89
rect 402 -90 403 -89
rect 403 -90 404 -89
rect 404 -90 405 -89
rect 405 -90 406 -89
rect 406 -90 407 -89
rect 407 -90 408 -89
rect 408 -90 409 -89
rect 409 -90 410 -89
rect 410 -90 411 -89
rect 411 -90 412 -89
rect 412 -90 413 -89
rect 413 -90 414 -89
rect 414 -90 415 -89
rect 415 -90 416 -89
rect 416 -90 417 -89
rect 417 -90 418 -89
rect 418 -90 419 -89
rect 419 -90 420 -89
rect 420 -90 421 -89
rect 421 -90 422 -89
rect 422 -90 423 -89
rect 423 -90 424 -89
rect 424 -90 425 -89
rect 425 -90 426 -89
rect 426 -90 427 -89
rect 427 -90 428 -89
rect 428 -90 429 -89
rect 429 -90 430 -89
rect 430 -90 431 -89
rect 431 -90 432 -89
rect 432 -90 433 -89
rect 433 -90 434 -89
rect 434 -90 435 -89
rect 435 -90 436 -89
rect 436 -90 437 -89
rect 437 -90 438 -89
rect 438 -90 439 -89
rect 439 -90 440 -89
rect 440 -90 441 -89
rect 441 -90 442 -89
rect 442 -90 443 -89
rect 443 -90 444 -89
rect 444 -90 445 -89
rect 445 -90 446 -89
rect 446 -90 447 -89
rect 447 -90 448 -89
rect 448 -90 449 -89
rect 449 -90 450 -89
rect 450 -90 451 -89
rect 451 -90 452 -89
rect 452 -90 453 -89
rect 453 -90 454 -89
rect 454 -90 455 -89
rect 455 -90 456 -89
rect 456 -90 457 -89
rect 457 -90 458 -89
rect 458 -90 459 -89
rect 459 -90 460 -89
rect 460 -90 461 -89
rect 461 -90 462 -89
rect 462 -90 463 -89
rect 463 -90 464 -89
rect 464 -90 465 -89
rect 465 -90 466 -89
rect 466 -90 467 -89
rect 467 -90 468 -89
rect 468 -90 469 -89
rect 469 -90 470 -89
rect 470 -90 471 -89
rect 471 -90 472 -89
rect 472 -90 473 -89
rect 473 -90 474 -89
rect 474 -90 475 -89
rect 475 -90 476 -89
rect 476 -90 477 -89
rect 477 -90 478 -89
rect 478 -90 479 -89
rect 479 -90 480 -89
rect 2 -91 3 -90
rect 3 -91 4 -90
rect 4 -91 5 -90
rect 5 -91 6 -90
rect 6 -91 7 -90
rect 7 -91 8 -90
rect 8 -91 9 -90
rect 9 -91 10 -90
rect 10 -91 11 -90
rect 11 -91 12 -90
rect 12 -91 13 -90
rect 13 -91 14 -90
rect 19 -91 20 -90
rect 20 -91 21 -90
rect 21 -91 22 -90
rect 22 -91 23 -90
rect 23 -91 24 -90
rect 24 -91 25 -90
rect 25 -91 26 -90
rect 26 -91 27 -90
rect 27 -91 28 -90
rect 28 -91 29 -90
rect 29 -91 30 -90
rect 30 -91 31 -90
rect 31 -91 32 -90
rect 32 -91 33 -90
rect 33 -91 34 -90
rect 34 -91 35 -90
rect 35 -91 36 -90
rect 36 -91 37 -90
rect 37 -91 38 -90
rect 38 -91 39 -90
rect 39 -91 40 -90
rect 40 -91 41 -90
rect 41 -91 42 -90
rect 42 -91 43 -90
rect 43 -91 44 -90
rect 44 -91 45 -90
rect 45 -91 46 -90
rect 51 -91 52 -90
rect 52 -91 53 -90
rect 53 -91 54 -90
rect 54 -91 55 -90
rect 55 -91 56 -90
rect 56 -91 57 -90
rect 57 -91 58 -90
rect 58 -91 59 -90
rect 59 -91 60 -90
rect 60 -91 61 -90
rect 61 -91 62 -90
rect 62 -91 63 -90
rect 63 -91 64 -90
rect 64 -91 65 -90
rect 65 -91 66 -90
rect 66 -91 67 -90
rect 67 -91 68 -90
rect 68 -91 69 -90
rect 69 -91 70 -90
rect 70 -91 71 -90
rect 71 -91 72 -90
rect 72 -91 73 -90
rect 73 -91 74 -90
rect 74 -91 75 -90
rect 75 -91 76 -90
rect 76 -91 77 -90
rect 77 -91 78 -90
rect 83 -91 84 -90
rect 84 -91 85 -90
rect 85 -91 86 -90
rect 86 -91 87 -90
rect 87 -91 88 -90
rect 88 -91 89 -90
rect 89 -91 90 -90
rect 90 -91 91 -90
rect 91 -91 92 -90
rect 92 -91 93 -90
rect 93 -91 94 -90
rect 94 -91 95 -90
rect 95 -91 96 -90
rect 96 -91 97 -90
rect 97 -91 98 -90
rect 98 -91 99 -90
rect 99 -91 100 -90
rect 100 -91 101 -90
rect 101 -91 102 -90
rect 102 -91 103 -90
rect 103 -91 104 -90
rect 104 -91 105 -90
rect 105 -91 106 -90
rect 106 -91 107 -90
rect 107 -91 108 -90
rect 108 -91 109 -90
rect 109 -91 110 -90
rect 115 -91 116 -90
rect 116 -91 117 -90
rect 117 -91 118 -90
rect 118 -91 119 -90
rect 119 -91 120 -90
rect 120 -91 121 -90
rect 121 -91 122 -90
rect 122 -91 123 -90
rect 123 -91 124 -90
rect 124 -91 125 -90
rect 125 -91 126 -90
rect 126 -91 127 -90
rect 127 -91 128 -90
rect 128 -91 129 -90
rect 129 -91 130 -90
rect 130 -91 131 -90
rect 131 -91 132 -90
rect 132 -91 133 -90
rect 133 -91 134 -90
rect 134 -91 135 -90
rect 135 -91 136 -90
rect 136 -91 137 -90
rect 137 -91 138 -90
rect 138 -91 139 -90
rect 139 -91 140 -90
rect 140 -91 141 -90
rect 141 -91 142 -90
rect 147 -91 148 -90
rect 148 -91 149 -90
rect 149 -91 150 -90
rect 150 -91 151 -90
rect 151 -91 152 -90
rect 152 -91 153 -90
rect 153 -91 154 -90
rect 154 -91 155 -90
rect 155 -91 156 -90
rect 156 -91 157 -90
rect 157 -91 158 -90
rect 158 -91 159 -90
rect 159 -91 160 -90
rect 160 -91 161 -90
rect 161 -91 162 -90
rect 162 -91 163 -90
rect 163 -91 164 -90
rect 164 -91 165 -90
rect 165 -91 166 -90
rect 166 -91 167 -90
rect 167 -91 168 -90
rect 168 -91 169 -90
rect 169 -91 170 -90
rect 170 -91 171 -90
rect 171 -91 172 -90
rect 172 -91 173 -90
rect 173 -91 174 -90
rect 179 -91 180 -90
rect 180 -91 181 -90
rect 181 -91 182 -90
rect 182 -91 183 -90
rect 183 -91 184 -90
rect 184 -91 185 -90
rect 185 -91 186 -90
rect 186 -91 187 -90
rect 187 -91 188 -90
rect 188 -91 189 -90
rect 189 -91 190 -90
rect 190 -91 191 -90
rect 191 -91 192 -90
rect 192 -91 193 -90
rect 193 -91 194 -90
rect 194 -91 195 -90
rect 195 -91 196 -90
rect 196 -91 197 -90
rect 197 -91 198 -90
rect 198 -91 199 -90
rect 199 -91 200 -90
rect 200 -91 201 -90
rect 201 -91 202 -90
rect 202 -91 203 -90
rect 203 -91 204 -90
rect 204 -91 205 -90
rect 205 -91 206 -90
rect 206 -91 207 -90
rect 207 -91 208 -90
rect 208 -91 209 -90
rect 209 -91 210 -90
rect 210 -91 211 -90
rect 211 -91 212 -90
rect 212 -91 213 -90
rect 213 -91 214 -90
rect 214 -91 215 -90
rect 215 -91 216 -90
rect 216 -91 217 -90
rect 217 -91 218 -90
rect 218 -91 219 -90
rect 219 -91 220 -90
rect 220 -91 221 -90
rect 221 -91 222 -90
rect 222 -91 223 -90
rect 223 -91 224 -90
rect 224 -91 225 -90
rect 225 -91 226 -90
rect 226 -91 227 -90
rect 227 -91 228 -90
rect 228 -91 229 -90
rect 229 -91 230 -90
rect 230 -91 231 -90
rect 231 -91 232 -90
rect 232 -91 233 -90
rect 233 -91 234 -90
rect 234 -91 235 -90
rect 235 -91 236 -90
rect 236 -91 237 -90
rect 237 -91 238 -90
rect 238 -91 239 -90
rect 239 -91 240 -90
rect 240 -91 241 -90
rect 241 -91 242 -90
rect 242 -91 243 -90
rect 243 -91 244 -90
rect 244 -91 245 -90
rect 245 -91 246 -90
rect 246 -91 247 -90
rect 247 -91 248 -90
rect 248 -91 249 -90
rect 249 -91 250 -90
rect 250 -91 251 -90
rect 251 -91 252 -90
rect 252 -91 253 -90
rect 253 -91 254 -90
rect 254 -91 255 -90
rect 255 -91 256 -90
rect 256 -91 257 -90
rect 257 -91 258 -90
rect 258 -91 259 -90
rect 259 -91 260 -90
rect 260 -91 261 -90
rect 261 -91 262 -90
rect 262 -91 263 -90
rect 263 -91 264 -90
rect 264 -91 265 -90
rect 265 -91 266 -90
rect 266 -91 267 -90
rect 267 -91 268 -90
rect 268 -91 269 -90
rect 269 -91 270 -90
rect 270 -91 271 -90
rect 271 -91 272 -90
rect 272 -91 273 -90
rect 273 -91 274 -90
rect 274 -91 275 -90
rect 275 -91 276 -90
rect 276 -91 277 -90
rect 277 -91 278 -90
rect 278 -91 279 -90
rect 279 -91 280 -90
rect 280 -91 281 -90
rect 281 -91 282 -90
rect 282 -91 283 -90
rect 283 -91 284 -90
rect 284 -91 285 -90
rect 285 -91 286 -90
rect 286 -91 287 -90
rect 287 -91 288 -90
rect 288 -91 289 -90
rect 289 -91 290 -90
rect 290 -91 291 -90
rect 291 -91 292 -90
rect 292 -91 293 -90
rect 293 -91 294 -90
rect 294 -91 295 -90
rect 295 -91 296 -90
rect 296 -91 297 -90
rect 297 -91 298 -90
rect 298 -91 299 -90
rect 299 -91 300 -90
rect 300 -91 301 -90
rect 301 -91 302 -90
rect 302 -91 303 -90
rect 303 -91 304 -90
rect 304 -91 305 -90
rect 305 -91 306 -90
rect 306 -91 307 -90
rect 307 -91 308 -90
rect 308 -91 309 -90
rect 309 -91 310 -90
rect 310 -91 311 -90
rect 311 -91 312 -90
rect 312 -91 313 -90
rect 313 -91 314 -90
rect 314 -91 315 -90
rect 315 -91 316 -90
rect 316 -91 317 -90
rect 317 -91 318 -90
rect 318 -91 319 -90
rect 319 -91 320 -90
rect 320 -91 321 -90
rect 321 -91 322 -90
rect 322 -91 323 -90
rect 323 -91 324 -90
rect 324 -91 325 -90
rect 325 -91 326 -90
rect 326 -91 327 -90
rect 327 -91 328 -90
rect 328 -91 329 -90
rect 329 -91 330 -90
rect 330 -91 331 -90
rect 331 -91 332 -90
rect 332 -91 333 -90
rect 333 -91 334 -90
rect 334 -91 335 -90
rect 335 -91 336 -90
rect 336 -91 337 -90
rect 337 -91 338 -90
rect 338 -91 339 -90
rect 339 -91 340 -90
rect 340 -91 341 -90
rect 341 -91 342 -90
rect 342 -91 343 -90
rect 343 -91 344 -90
rect 344 -91 345 -90
rect 345 -91 346 -90
rect 346 -91 347 -90
rect 347 -91 348 -90
rect 348 -91 349 -90
rect 349 -91 350 -90
rect 350 -91 351 -90
rect 351 -91 352 -90
rect 352 -91 353 -90
rect 353 -91 354 -90
rect 354 -91 355 -90
rect 355 -91 356 -90
rect 356 -91 357 -90
rect 357 -91 358 -90
rect 358 -91 359 -90
rect 359 -91 360 -90
rect 360 -91 361 -90
rect 361 -91 362 -90
rect 362 -91 363 -90
rect 363 -91 364 -90
rect 364 -91 365 -90
rect 365 -91 366 -90
rect 366 -91 367 -90
rect 367 -91 368 -90
rect 368 -91 369 -90
rect 369 -91 370 -90
rect 370 -91 371 -90
rect 371 -91 372 -90
rect 372 -91 373 -90
rect 373 -91 374 -90
rect 374 -91 375 -90
rect 375 -91 376 -90
rect 376 -91 377 -90
rect 377 -91 378 -90
rect 378 -91 379 -90
rect 379 -91 380 -90
rect 380 -91 381 -90
rect 381 -91 382 -90
rect 382 -91 383 -90
rect 383 -91 384 -90
rect 384 -91 385 -90
rect 385 -91 386 -90
rect 386 -91 387 -90
rect 387 -91 388 -90
rect 388 -91 389 -90
rect 389 -91 390 -90
rect 390 -91 391 -90
rect 391 -91 392 -90
rect 392 -91 393 -90
rect 393 -91 394 -90
rect 394 -91 395 -90
rect 395 -91 396 -90
rect 396 -91 397 -90
rect 397 -91 398 -90
rect 398 -91 399 -90
rect 399 -91 400 -90
rect 400 -91 401 -90
rect 401 -91 402 -90
rect 402 -91 403 -90
rect 403 -91 404 -90
rect 404 -91 405 -90
rect 405 -91 406 -90
rect 406 -91 407 -90
rect 407 -91 408 -90
rect 408 -91 409 -90
rect 409 -91 410 -90
rect 410 -91 411 -90
rect 411 -91 412 -90
rect 412 -91 413 -90
rect 413 -91 414 -90
rect 414 -91 415 -90
rect 415 -91 416 -90
rect 416 -91 417 -90
rect 417 -91 418 -90
rect 418 -91 419 -90
rect 419 -91 420 -90
rect 420 -91 421 -90
rect 421 -91 422 -90
rect 422 -91 423 -90
rect 423 -91 424 -90
rect 424 -91 425 -90
rect 425 -91 426 -90
rect 426 -91 427 -90
rect 427 -91 428 -90
rect 428 -91 429 -90
rect 429 -91 430 -90
rect 430 -91 431 -90
rect 431 -91 432 -90
rect 432 -91 433 -90
rect 433 -91 434 -90
rect 434 -91 435 -90
rect 435 -91 436 -90
rect 436 -91 437 -90
rect 437 -91 438 -90
rect 438 -91 439 -90
rect 439 -91 440 -90
rect 440 -91 441 -90
rect 441 -91 442 -90
rect 442 -91 443 -90
rect 443 -91 444 -90
rect 444 -91 445 -90
rect 445 -91 446 -90
rect 446 -91 447 -90
rect 447 -91 448 -90
rect 448 -91 449 -90
rect 449 -91 450 -90
rect 450 -91 451 -90
rect 451 -91 452 -90
rect 452 -91 453 -90
rect 453 -91 454 -90
rect 454 -91 455 -90
rect 455 -91 456 -90
rect 456 -91 457 -90
rect 457 -91 458 -90
rect 458 -91 459 -90
rect 459 -91 460 -90
rect 460 -91 461 -90
rect 461 -91 462 -90
rect 462 -91 463 -90
rect 463 -91 464 -90
rect 464 -91 465 -90
rect 465 -91 466 -90
rect 466 -91 467 -90
rect 467 -91 468 -90
rect 468 -91 469 -90
rect 469 -91 470 -90
rect 470 -91 471 -90
rect 471 -91 472 -90
rect 472 -91 473 -90
rect 473 -91 474 -90
rect 474 -91 475 -90
rect 475 -91 476 -90
rect 476 -91 477 -90
rect 477 -91 478 -90
rect 478 -91 479 -90
rect 479 -91 480 -90
rect 2 -92 3 -91
rect 3 -92 4 -91
rect 4 -92 5 -91
rect 5 -92 6 -91
rect 6 -92 7 -91
rect 7 -92 8 -91
rect 25 -92 26 -91
rect 26 -92 27 -91
rect 27 -92 28 -91
rect 28 -92 29 -91
rect 29 -92 30 -91
rect 30 -92 31 -91
rect 31 -92 32 -91
rect 32 -92 33 -91
rect 33 -92 34 -91
rect 34 -92 35 -91
rect 35 -92 36 -91
rect 36 -92 37 -91
rect 37 -92 38 -91
rect 38 -92 39 -91
rect 39 -92 40 -91
rect 57 -92 58 -91
rect 58 -92 59 -91
rect 59 -92 60 -91
rect 60 -92 61 -91
rect 61 -92 62 -91
rect 62 -92 63 -91
rect 63 -92 64 -91
rect 64 -92 65 -91
rect 65 -92 66 -91
rect 66 -92 67 -91
rect 67 -92 68 -91
rect 68 -92 69 -91
rect 69 -92 70 -91
rect 70 -92 71 -91
rect 71 -92 72 -91
rect 89 -92 90 -91
rect 90 -92 91 -91
rect 91 -92 92 -91
rect 92 -92 93 -91
rect 93 -92 94 -91
rect 94 -92 95 -91
rect 95 -92 96 -91
rect 96 -92 97 -91
rect 97 -92 98 -91
rect 98 -92 99 -91
rect 99 -92 100 -91
rect 100 -92 101 -91
rect 101 -92 102 -91
rect 102 -92 103 -91
rect 103 -92 104 -91
rect 121 -92 122 -91
rect 122 -92 123 -91
rect 123 -92 124 -91
rect 124 -92 125 -91
rect 125 -92 126 -91
rect 126 -92 127 -91
rect 127 -92 128 -91
rect 128 -92 129 -91
rect 129 -92 130 -91
rect 130 -92 131 -91
rect 131 -92 132 -91
rect 132 -92 133 -91
rect 133 -92 134 -91
rect 134 -92 135 -91
rect 135 -92 136 -91
rect 153 -92 154 -91
rect 154 -92 155 -91
rect 155 -92 156 -91
rect 156 -92 157 -91
rect 157 -92 158 -91
rect 158 -92 159 -91
rect 159 -92 160 -91
rect 160 -92 161 -91
rect 161 -92 162 -91
rect 162 -92 163 -91
rect 163 -92 164 -91
rect 164 -92 165 -91
rect 165 -92 166 -91
rect 166 -92 167 -91
rect 167 -92 168 -91
rect 185 -92 186 -91
rect 186 -92 187 -91
rect 187 -92 188 -91
rect 188 -92 189 -91
rect 189 -92 190 -91
rect 190 -92 191 -91
rect 191 -92 192 -91
rect 192 -92 193 -91
rect 193 -92 194 -91
rect 194 -92 195 -91
rect 195 -92 196 -91
rect 196 -92 197 -91
rect 197 -92 198 -91
rect 198 -92 199 -91
rect 199 -92 200 -91
rect 200 -92 201 -91
rect 201 -92 202 -91
rect 202 -92 203 -91
rect 203 -92 204 -91
rect 204 -92 205 -91
rect 205 -92 206 -91
rect 206 -92 207 -91
rect 207 -92 208 -91
rect 208 -92 209 -91
rect 209 -92 210 -91
rect 210 -92 211 -91
rect 211 -92 212 -91
rect 212 -92 213 -91
rect 213 -92 214 -91
rect 214 -92 215 -91
rect 215 -92 216 -91
rect 216 -92 217 -91
rect 217 -92 218 -91
rect 218 -92 219 -91
rect 219 -92 220 -91
rect 220 -92 221 -91
rect 221 -92 222 -91
rect 222 -92 223 -91
rect 223 -92 224 -91
rect 224 -92 225 -91
rect 225 -92 226 -91
rect 226 -92 227 -91
rect 227 -92 228 -91
rect 228 -92 229 -91
rect 229 -92 230 -91
rect 230 -92 231 -91
rect 231 -92 232 -91
rect 232 -92 233 -91
rect 233 -92 234 -91
rect 234 -92 235 -91
rect 235 -92 236 -91
rect 236 -92 237 -91
rect 237 -92 238 -91
rect 238 -92 239 -91
rect 239 -92 240 -91
rect 240 -92 241 -91
rect 241 -92 242 -91
rect 242 -92 243 -91
rect 243 -92 244 -91
rect 244 -92 245 -91
rect 245 -92 246 -91
rect 246 -92 247 -91
rect 247 -92 248 -91
rect 248 -92 249 -91
rect 249 -92 250 -91
rect 250 -92 251 -91
rect 251 -92 252 -91
rect 252 -92 253 -91
rect 253 -92 254 -91
rect 254 -92 255 -91
rect 255 -92 256 -91
rect 256 -92 257 -91
rect 257 -92 258 -91
rect 258 -92 259 -91
rect 259 -92 260 -91
rect 260 -92 261 -91
rect 261 -92 262 -91
rect 262 -92 263 -91
rect 263 -92 264 -91
rect 264 -92 265 -91
rect 265 -92 266 -91
rect 266 -92 267 -91
rect 267 -92 268 -91
rect 268 -92 269 -91
rect 269 -92 270 -91
rect 270 -92 271 -91
rect 271 -92 272 -91
rect 272 -92 273 -91
rect 273 -92 274 -91
rect 274 -92 275 -91
rect 275 -92 276 -91
rect 276 -92 277 -91
rect 277 -92 278 -91
rect 278 -92 279 -91
rect 279 -92 280 -91
rect 280 -92 281 -91
rect 281 -92 282 -91
rect 282 -92 283 -91
rect 283 -92 284 -91
rect 284 -92 285 -91
rect 285 -92 286 -91
rect 286 -92 287 -91
rect 287 -92 288 -91
rect 288 -92 289 -91
rect 289 -92 290 -91
rect 290 -92 291 -91
rect 291 -92 292 -91
rect 292 -92 293 -91
rect 293 -92 294 -91
rect 294 -92 295 -91
rect 295 -92 296 -91
rect 296 -92 297 -91
rect 297 -92 298 -91
rect 298 -92 299 -91
rect 299 -92 300 -91
rect 300 -92 301 -91
rect 301 -92 302 -91
rect 302 -92 303 -91
rect 303 -92 304 -91
rect 304 -92 305 -91
rect 305 -92 306 -91
rect 306 -92 307 -91
rect 307 -92 308 -91
rect 308 -92 309 -91
rect 309 -92 310 -91
rect 310 -92 311 -91
rect 311 -92 312 -91
rect 312 -92 313 -91
rect 313 -92 314 -91
rect 314 -92 315 -91
rect 315 -92 316 -91
rect 316 -92 317 -91
rect 317 -92 318 -91
rect 318 -92 319 -91
rect 319 -92 320 -91
rect 320 -92 321 -91
rect 321 -92 322 -91
rect 322 -92 323 -91
rect 323 -92 324 -91
rect 324 -92 325 -91
rect 325 -92 326 -91
rect 326 -92 327 -91
rect 327 -92 328 -91
rect 328 -92 329 -91
rect 329 -92 330 -91
rect 330 -92 331 -91
rect 331 -92 332 -91
rect 332 -92 333 -91
rect 333 -92 334 -91
rect 334 -92 335 -91
rect 335 -92 336 -91
rect 336 -92 337 -91
rect 337 -92 338 -91
rect 338 -92 339 -91
rect 339 -92 340 -91
rect 340 -92 341 -91
rect 341 -92 342 -91
rect 342 -92 343 -91
rect 343 -92 344 -91
rect 344 -92 345 -91
rect 345 -92 346 -91
rect 346 -92 347 -91
rect 347 -92 348 -91
rect 348 -92 349 -91
rect 349 -92 350 -91
rect 350 -92 351 -91
rect 351 -92 352 -91
rect 352 -92 353 -91
rect 353 -92 354 -91
rect 354 -92 355 -91
rect 355 -92 356 -91
rect 356 -92 357 -91
rect 357 -92 358 -91
rect 358 -92 359 -91
rect 359 -92 360 -91
rect 360 -92 361 -91
rect 361 -92 362 -91
rect 362 -92 363 -91
rect 363 -92 364 -91
rect 364 -92 365 -91
rect 365 -92 366 -91
rect 366 -92 367 -91
rect 367 -92 368 -91
rect 368 -92 369 -91
rect 369 -92 370 -91
rect 370 -92 371 -91
rect 371 -92 372 -91
rect 372 -92 373 -91
rect 373 -92 374 -91
rect 374 -92 375 -91
rect 375 -92 376 -91
rect 376 -92 377 -91
rect 377 -92 378 -91
rect 378 -92 379 -91
rect 379 -92 380 -91
rect 380 -92 381 -91
rect 381 -92 382 -91
rect 382 -92 383 -91
rect 383 -92 384 -91
rect 384 -92 385 -91
rect 385 -92 386 -91
rect 386 -92 387 -91
rect 387 -92 388 -91
rect 388 -92 389 -91
rect 389 -92 390 -91
rect 390 -92 391 -91
rect 391 -92 392 -91
rect 392 -92 393 -91
rect 393 -92 394 -91
rect 394 -92 395 -91
rect 395 -92 396 -91
rect 396 -92 397 -91
rect 397 -92 398 -91
rect 398 -92 399 -91
rect 399 -92 400 -91
rect 400 -92 401 -91
rect 401 -92 402 -91
rect 402 -92 403 -91
rect 403 -92 404 -91
rect 404 -92 405 -91
rect 405 -92 406 -91
rect 406 -92 407 -91
rect 407 -92 408 -91
rect 408 -92 409 -91
rect 409 -92 410 -91
rect 410 -92 411 -91
rect 411 -92 412 -91
rect 412 -92 413 -91
rect 413 -92 414 -91
rect 414 -92 415 -91
rect 415 -92 416 -91
rect 416 -92 417 -91
rect 417 -92 418 -91
rect 418 -92 419 -91
rect 419 -92 420 -91
rect 420 -92 421 -91
rect 421 -92 422 -91
rect 422 -92 423 -91
rect 423 -92 424 -91
rect 424 -92 425 -91
rect 425 -92 426 -91
rect 426 -92 427 -91
rect 427 -92 428 -91
rect 428 -92 429 -91
rect 429 -92 430 -91
rect 430 -92 431 -91
rect 431 -92 432 -91
rect 432 -92 433 -91
rect 433 -92 434 -91
rect 434 -92 435 -91
rect 435 -92 436 -91
rect 436 -92 437 -91
rect 437 -92 438 -91
rect 438 -92 439 -91
rect 439 -92 440 -91
rect 440 -92 441 -91
rect 441 -92 442 -91
rect 442 -92 443 -91
rect 443 -92 444 -91
rect 444 -92 445 -91
rect 445 -92 446 -91
rect 446 -92 447 -91
rect 447 -92 448 -91
rect 448 -92 449 -91
rect 449 -92 450 -91
rect 450 -92 451 -91
rect 451 -92 452 -91
rect 452 -92 453 -91
rect 453 -92 454 -91
rect 454 -92 455 -91
rect 455 -92 456 -91
rect 456 -92 457 -91
rect 457 -92 458 -91
rect 458 -92 459 -91
rect 459 -92 460 -91
rect 460 -92 461 -91
rect 461 -92 462 -91
rect 462 -92 463 -91
rect 463 -92 464 -91
rect 464 -92 465 -91
rect 465 -92 466 -91
rect 466 -92 467 -91
rect 467 -92 468 -91
rect 468 -92 469 -91
rect 469 -92 470 -91
rect 470 -92 471 -91
rect 471 -92 472 -91
rect 472 -92 473 -91
rect 473 -92 474 -91
rect 474 -92 475 -91
rect 475 -92 476 -91
rect 476 -92 477 -91
rect 477 -92 478 -91
rect 478 -92 479 -91
rect 479 -92 480 -91
rect 2 -93 3 -92
rect 3 -93 4 -92
rect 4 -93 5 -92
rect 5 -93 6 -92
rect 6 -93 7 -92
rect 7 -93 8 -92
rect 8 -93 9 -92
rect 25 -93 26 -92
rect 26 -93 27 -92
rect 27 -93 28 -92
rect 28 -93 29 -92
rect 29 -93 30 -92
rect 30 -93 31 -92
rect 31 -93 32 -92
rect 32 -93 33 -92
rect 33 -93 34 -92
rect 34 -93 35 -92
rect 35 -93 36 -92
rect 36 -93 37 -92
rect 37 -93 38 -92
rect 38 -93 39 -92
rect 39 -93 40 -92
rect 40 -93 41 -92
rect 57 -93 58 -92
rect 58 -93 59 -92
rect 59 -93 60 -92
rect 60 -93 61 -92
rect 61 -93 62 -92
rect 62 -93 63 -92
rect 63 -93 64 -92
rect 64 -93 65 -92
rect 65 -93 66 -92
rect 66 -93 67 -92
rect 67 -93 68 -92
rect 68 -93 69 -92
rect 69 -93 70 -92
rect 70 -93 71 -92
rect 71 -93 72 -92
rect 72 -93 73 -92
rect 89 -93 90 -92
rect 90 -93 91 -92
rect 91 -93 92 -92
rect 92 -93 93 -92
rect 93 -93 94 -92
rect 94 -93 95 -92
rect 95 -93 96 -92
rect 96 -93 97 -92
rect 97 -93 98 -92
rect 98 -93 99 -92
rect 99 -93 100 -92
rect 100 -93 101 -92
rect 101 -93 102 -92
rect 102 -93 103 -92
rect 103 -93 104 -92
rect 104 -93 105 -92
rect 121 -93 122 -92
rect 122 -93 123 -92
rect 123 -93 124 -92
rect 124 -93 125 -92
rect 125 -93 126 -92
rect 126 -93 127 -92
rect 127 -93 128 -92
rect 128 -93 129 -92
rect 129 -93 130 -92
rect 130 -93 131 -92
rect 131 -93 132 -92
rect 132 -93 133 -92
rect 133 -93 134 -92
rect 134 -93 135 -92
rect 135 -93 136 -92
rect 136 -93 137 -92
rect 153 -93 154 -92
rect 154 -93 155 -92
rect 155 -93 156 -92
rect 156 -93 157 -92
rect 157 -93 158 -92
rect 158 -93 159 -92
rect 159 -93 160 -92
rect 160 -93 161 -92
rect 161 -93 162 -92
rect 162 -93 163 -92
rect 163 -93 164 -92
rect 164 -93 165 -92
rect 165 -93 166 -92
rect 166 -93 167 -92
rect 167 -93 168 -92
rect 168 -93 169 -92
rect 185 -93 186 -92
rect 186 -93 187 -92
rect 187 -93 188 -92
rect 188 -93 189 -92
rect 189 -93 190 -92
rect 190 -93 191 -92
rect 191 -93 192 -92
rect 192 -93 193 -92
rect 193 -93 194 -92
rect 194 -93 195 -92
rect 195 -93 196 -92
rect 196 -93 197 -92
rect 197 -93 198 -92
rect 198 -93 199 -92
rect 199 -93 200 -92
rect 200 -93 201 -92
rect 201 -93 202 -92
rect 202 -93 203 -92
rect 203 -93 204 -92
rect 204 -93 205 -92
rect 205 -93 206 -92
rect 206 -93 207 -92
rect 207 -93 208 -92
rect 208 -93 209 -92
rect 209 -93 210 -92
rect 210 -93 211 -92
rect 211 -93 212 -92
rect 212 -93 213 -92
rect 213 -93 214 -92
rect 214 -93 215 -92
rect 215 -93 216 -92
rect 216 -93 217 -92
rect 217 -93 218 -92
rect 218 -93 219 -92
rect 219 -93 220 -92
rect 220 -93 221 -92
rect 221 -93 222 -92
rect 222 -93 223 -92
rect 223 -93 224 -92
rect 224 -93 225 -92
rect 225 -93 226 -92
rect 226 -93 227 -92
rect 227 -93 228 -92
rect 228 -93 229 -92
rect 229 -93 230 -92
rect 230 -93 231 -92
rect 231 -93 232 -92
rect 232 -93 233 -92
rect 233 -93 234 -92
rect 234 -93 235 -92
rect 235 -93 236 -92
rect 236 -93 237 -92
rect 237 -93 238 -92
rect 238 -93 239 -92
rect 239 -93 240 -92
rect 240 -93 241 -92
rect 241 -93 242 -92
rect 242 -93 243 -92
rect 243 -93 244 -92
rect 244 -93 245 -92
rect 245 -93 246 -92
rect 246 -93 247 -92
rect 247 -93 248 -92
rect 248 -93 249 -92
rect 249 -93 250 -92
rect 250 -93 251 -92
rect 251 -93 252 -92
rect 252 -93 253 -92
rect 253 -93 254 -92
rect 254 -93 255 -92
rect 255 -93 256 -92
rect 256 -93 257 -92
rect 257 -93 258 -92
rect 258 -93 259 -92
rect 259 -93 260 -92
rect 260 -93 261 -92
rect 261 -93 262 -92
rect 262 -93 263 -92
rect 263 -93 264 -92
rect 264 -93 265 -92
rect 265 -93 266 -92
rect 266 -93 267 -92
rect 267 -93 268 -92
rect 268 -93 269 -92
rect 269 -93 270 -92
rect 270 -93 271 -92
rect 271 -93 272 -92
rect 272 -93 273 -92
rect 273 -93 274 -92
rect 274 -93 275 -92
rect 275 -93 276 -92
rect 276 -93 277 -92
rect 277 -93 278 -92
rect 278 -93 279 -92
rect 279 -93 280 -92
rect 280 -93 281 -92
rect 281 -93 282 -92
rect 282 -93 283 -92
rect 283 -93 284 -92
rect 284 -93 285 -92
rect 285 -93 286 -92
rect 286 -93 287 -92
rect 287 -93 288 -92
rect 288 -93 289 -92
rect 289 -93 290 -92
rect 290 -93 291 -92
rect 291 -93 292 -92
rect 292 -93 293 -92
rect 293 -93 294 -92
rect 294 -93 295 -92
rect 295 -93 296 -92
rect 296 -93 297 -92
rect 297 -93 298 -92
rect 298 -93 299 -92
rect 299 -93 300 -92
rect 300 -93 301 -92
rect 301 -93 302 -92
rect 302 -93 303 -92
rect 303 -93 304 -92
rect 304 -93 305 -92
rect 305 -93 306 -92
rect 306 -93 307 -92
rect 307 -93 308 -92
rect 308 -93 309 -92
rect 309 -93 310 -92
rect 310 -93 311 -92
rect 311 -93 312 -92
rect 312 -93 313 -92
rect 313 -93 314 -92
rect 314 -93 315 -92
rect 315 -93 316 -92
rect 316 -93 317 -92
rect 317 -93 318 -92
rect 318 -93 319 -92
rect 319 -93 320 -92
rect 320 -93 321 -92
rect 321 -93 322 -92
rect 322 -93 323 -92
rect 323 -93 324 -92
rect 324 -93 325 -92
rect 325 -93 326 -92
rect 326 -93 327 -92
rect 327 -93 328 -92
rect 328 -93 329 -92
rect 329 -93 330 -92
rect 330 -93 331 -92
rect 331 -93 332 -92
rect 332 -93 333 -92
rect 333 -93 334 -92
rect 334 -93 335 -92
rect 335 -93 336 -92
rect 336 -93 337 -92
rect 337 -93 338 -92
rect 338 -93 339 -92
rect 339 -93 340 -92
rect 340 -93 341 -92
rect 341 -93 342 -92
rect 342 -93 343 -92
rect 343 -93 344 -92
rect 344 -93 345 -92
rect 345 -93 346 -92
rect 346 -93 347 -92
rect 347 -93 348 -92
rect 348 -93 349 -92
rect 349 -93 350 -92
rect 350 -93 351 -92
rect 351 -93 352 -92
rect 352 -93 353 -92
rect 353 -93 354 -92
rect 354 -93 355 -92
rect 355 -93 356 -92
rect 356 -93 357 -92
rect 357 -93 358 -92
rect 358 -93 359 -92
rect 359 -93 360 -92
rect 360 -93 361 -92
rect 361 -93 362 -92
rect 362 -93 363 -92
rect 363 -93 364 -92
rect 364 -93 365 -92
rect 365 -93 366 -92
rect 366 -93 367 -92
rect 367 -93 368 -92
rect 368 -93 369 -92
rect 369 -93 370 -92
rect 370 -93 371 -92
rect 371 -93 372 -92
rect 372 -93 373 -92
rect 373 -93 374 -92
rect 374 -93 375 -92
rect 375 -93 376 -92
rect 376 -93 377 -92
rect 377 -93 378 -92
rect 378 -93 379 -92
rect 379 -93 380 -92
rect 380 -93 381 -92
rect 381 -93 382 -92
rect 382 -93 383 -92
rect 383 -93 384 -92
rect 384 -93 385 -92
rect 385 -93 386 -92
rect 386 -93 387 -92
rect 387 -93 388 -92
rect 388 -93 389 -92
rect 389 -93 390 -92
rect 390 -93 391 -92
rect 391 -93 392 -92
rect 392 -93 393 -92
rect 393 -93 394 -92
rect 394 -93 395 -92
rect 395 -93 396 -92
rect 396 -93 397 -92
rect 397 -93 398 -92
rect 398 -93 399 -92
rect 399 -93 400 -92
rect 400 -93 401 -92
rect 401 -93 402 -92
rect 402 -93 403 -92
rect 403 -93 404 -92
rect 404 -93 405 -92
rect 405 -93 406 -92
rect 406 -93 407 -92
rect 407 -93 408 -92
rect 408 -93 409 -92
rect 409 -93 410 -92
rect 410 -93 411 -92
rect 411 -93 412 -92
rect 412 -93 413 -92
rect 413 -93 414 -92
rect 414 -93 415 -92
rect 415 -93 416 -92
rect 416 -93 417 -92
rect 417 -93 418 -92
rect 418 -93 419 -92
rect 419 -93 420 -92
rect 420 -93 421 -92
rect 421 -93 422 -92
rect 422 -93 423 -92
rect 423 -93 424 -92
rect 424 -93 425 -92
rect 425 -93 426 -92
rect 426 -93 427 -92
rect 427 -93 428 -92
rect 428 -93 429 -92
rect 429 -93 430 -92
rect 430 -93 431 -92
rect 431 -93 432 -92
rect 432 -93 433 -92
rect 433 -93 434 -92
rect 434 -93 435 -92
rect 435 -93 436 -92
rect 436 -93 437 -92
rect 437 -93 438 -92
rect 438 -93 439 -92
rect 439 -93 440 -92
rect 440 -93 441 -92
rect 441 -93 442 -92
rect 442 -93 443 -92
rect 443 -93 444 -92
rect 444 -93 445 -92
rect 445 -93 446 -92
rect 446 -93 447 -92
rect 447 -93 448 -92
rect 448 -93 449 -92
rect 449 -93 450 -92
rect 450 -93 451 -92
rect 451 -93 452 -92
rect 452 -93 453 -92
rect 453 -93 454 -92
rect 454 -93 455 -92
rect 455 -93 456 -92
rect 456 -93 457 -92
rect 457 -93 458 -92
rect 458 -93 459 -92
rect 459 -93 460 -92
rect 460 -93 461 -92
rect 461 -93 462 -92
rect 462 -93 463 -92
rect 463 -93 464 -92
rect 464 -93 465 -92
rect 465 -93 466 -92
rect 466 -93 467 -92
rect 467 -93 468 -92
rect 468 -93 469 -92
rect 469 -93 470 -92
rect 470 -93 471 -92
rect 471 -93 472 -92
rect 472 -93 473 -92
rect 473 -93 474 -92
rect 474 -93 475 -92
rect 475 -93 476 -92
rect 476 -93 477 -92
rect 477 -93 478 -92
rect 478 -93 479 -92
rect 479 -93 480 -92
rect 2 -94 3 -93
rect 3 -94 4 -93
rect 4 -94 5 -93
rect 5 -94 6 -93
rect 6 -94 7 -93
rect 7 -94 8 -93
rect 8 -94 9 -93
rect 9 -94 10 -93
rect 24 -94 25 -93
rect 25 -94 26 -93
rect 26 -94 27 -93
rect 27 -94 28 -93
rect 28 -94 29 -93
rect 29 -94 30 -93
rect 30 -94 31 -93
rect 31 -94 32 -93
rect 32 -94 33 -93
rect 33 -94 34 -93
rect 34 -94 35 -93
rect 35 -94 36 -93
rect 36 -94 37 -93
rect 37 -94 38 -93
rect 38 -94 39 -93
rect 39 -94 40 -93
rect 40 -94 41 -93
rect 41 -94 42 -93
rect 56 -94 57 -93
rect 57 -94 58 -93
rect 58 -94 59 -93
rect 59 -94 60 -93
rect 60 -94 61 -93
rect 61 -94 62 -93
rect 62 -94 63 -93
rect 63 -94 64 -93
rect 64 -94 65 -93
rect 65 -94 66 -93
rect 66 -94 67 -93
rect 67 -94 68 -93
rect 68 -94 69 -93
rect 69 -94 70 -93
rect 70 -94 71 -93
rect 71 -94 72 -93
rect 72 -94 73 -93
rect 88 -94 89 -93
rect 89 -94 90 -93
rect 90 -94 91 -93
rect 91 -94 92 -93
rect 92 -94 93 -93
rect 93 -94 94 -93
rect 94 -94 95 -93
rect 95 -94 96 -93
rect 96 -94 97 -93
rect 97 -94 98 -93
rect 98 -94 99 -93
rect 99 -94 100 -93
rect 100 -94 101 -93
rect 101 -94 102 -93
rect 102 -94 103 -93
rect 103 -94 104 -93
rect 104 -94 105 -93
rect 105 -94 106 -93
rect 120 -94 121 -93
rect 121 -94 122 -93
rect 122 -94 123 -93
rect 123 -94 124 -93
rect 124 -94 125 -93
rect 125 -94 126 -93
rect 126 -94 127 -93
rect 127 -94 128 -93
rect 128 -94 129 -93
rect 129 -94 130 -93
rect 130 -94 131 -93
rect 131 -94 132 -93
rect 132 -94 133 -93
rect 133 -94 134 -93
rect 134 -94 135 -93
rect 135 -94 136 -93
rect 136 -94 137 -93
rect 152 -94 153 -93
rect 153 -94 154 -93
rect 154 -94 155 -93
rect 155 -94 156 -93
rect 156 -94 157 -93
rect 157 -94 158 -93
rect 158 -94 159 -93
rect 159 -94 160 -93
rect 160 -94 161 -93
rect 161 -94 162 -93
rect 162 -94 163 -93
rect 163 -94 164 -93
rect 164 -94 165 -93
rect 165 -94 166 -93
rect 166 -94 167 -93
rect 167 -94 168 -93
rect 168 -94 169 -93
rect 169 -94 170 -93
rect 184 -94 185 -93
rect 185 -94 186 -93
rect 186 -94 187 -93
rect 187 -94 188 -93
rect 188 -94 189 -93
rect 189 -94 190 -93
rect 190 -94 191 -93
rect 191 -94 192 -93
rect 192 -94 193 -93
rect 193 -94 194 -93
rect 194 -94 195 -93
rect 195 -94 196 -93
rect 196 -94 197 -93
rect 197 -94 198 -93
rect 198 -94 199 -93
rect 199 -94 200 -93
rect 200 -94 201 -93
rect 201 -94 202 -93
rect 202 -94 203 -93
rect 203 -94 204 -93
rect 204 -94 205 -93
rect 205 -94 206 -93
rect 206 -94 207 -93
rect 207 -94 208 -93
rect 208 -94 209 -93
rect 209 -94 210 -93
rect 210 -94 211 -93
rect 211 -94 212 -93
rect 212 -94 213 -93
rect 213 -94 214 -93
rect 214 -94 215 -93
rect 215 -94 216 -93
rect 216 -94 217 -93
rect 217 -94 218 -93
rect 218 -94 219 -93
rect 219 -94 220 -93
rect 220 -94 221 -93
rect 221 -94 222 -93
rect 222 -94 223 -93
rect 223 -94 224 -93
rect 224 -94 225 -93
rect 225 -94 226 -93
rect 226 -94 227 -93
rect 227 -94 228 -93
rect 228 -94 229 -93
rect 229 -94 230 -93
rect 230 -94 231 -93
rect 231 -94 232 -93
rect 232 -94 233 -93
rect 233 -94 234 -93
rect 234 -94 235 -93
rect 235 -94 236 -93
rect 236 -94 237 -93
rect 237 -94 238 -93
rect 238 -94 239 -93
rect 239 -94 240 -93
rect 240 -94 241 -93
rect 241 -94 242 -93
rect 242 -94 243 -93
rect 243 -94 244 -93
rect 244 -94 245 -93
rect 245 -94 246 -93
rect 246 -94 247 -93
rect 247 -94 248 -93
rect 248 -94 249 -93
rect 249 -94 250 -93
rect 250 -94 251 -93
rect 251 -94 252 -93
rect 252 -94 253 -93
rect 253 -94 254 -93
rect 254 -94 255 -93
rect 255 -94 256 -93
rect 256 -94 257 -93
rect 257 -94 258 -93
rect 258 -94 259 -93
rect 259 -94 260 -93
rect 260 -94 261 -93
rect 261 -94 262 -93
rect 262 -94 263 -93
rect 263 -94 264 -93
rect 264 -94 265 -93
rect 265 -94 266 -93
rect 266 -94 267 -93
rect 267 -94 268 -93
rect 268 -94 269 -93
rect 269 -94 270 -93
rect 270 -94 271 -93
rect 271 -94 272 -93
rect 272 -94 273 -93
rect 273 -94 274 -93
rect 274 -94 275 -93
rect 275 -94 276 -93
rect 276 -94 277 -93
rect 277 -94 278 -93
rect 278 -94 279 -93
rect 279 -94 280 -93
rect 280 -94 281 -93
rect 281 -94 282 -93
rect 282 -94 283 -93
rect 283 -94 284 -93
rect 284 -94 285 -93
rect 285 -94 286 -93
rect 286 -94 287 -93
rect 287 -94 288 -93
rect 288 -94 289 -93
rect 289 -94 290 -93
rect 290 -94 291 -93
rect 291 -94 292 -93
rect 292 -94 293 -93
rect 293 -94 294 -93
rect 294 -94 295 -93
rect 295 -94 296 -93
rect 296 -94 297 -93
rect 297 -94 298 -93
rect 298 -94 299 -93
rect 299 -94 300 -93
rect 300 -94 301 -93
rect 301 -94 302 -93
rect 302 -94 303 -93
rect 303 -94 304 -93
rect 304 -94 305 -93
rect 305 -94 306 -93
rect 306 -94 307 -93
rect 307 -94 308 -93
rect 308 -94 309 -93
rect 309 -94 310 -93
rect 310 -94 311 -93
rect 311 -94 312 -93
rect 312 -94 313 -93
rect 313 -94 314 -93
rect 314 -94 315 -93
rect 315 -94 316 -93
rect 316 -94 317 -93
rect 317 -94 318 -93
rect 318 -94 319 -93
rect 319 -94 320 -93
rect 320 -94 321 -93
rect 321 -94 322 -93
rect 322 -94 323 -93
rect 323 -94 324 -93
rect 324 -94 325 -93
rect 325 -94 326 -93
rect 326 -94 327 -93
rect 327 -94 328 -93
rect 328 -94 329 -93
rect 329 -94 330 -93
rect 330 -94 331 -93
rect 331 -94 332 -93
rect 332 -94 333 -93
rect 333 -94 334 -93
rect 334 -94 335 -93
rect 335 -94 336 -93
rect 336 -94 337 -93
rect 337 -94 338 -93
rect 338 -94 339 -93
rect 339 -94 340 -93
rect 340 -94 341 -93
rect 341 -94 342 -93
rect 342 -94 343 -93
rect 343 -94 344 -93
rect 344 -94 345 -93
rect 345 -94 346 -93
rect 346 -94 347 -93
rect 347 -94 348 -93
rect 348 -94 349 -93
rect 349 -94 350 -93
rect 350 -94 351 -93
rect 351 -94 352 -93
rect 352 -94 353 -93
rect 353 -94 354 -93
rect 354 -94 355 -93
rect 355 -94 356 -93
rect 356 -94 357 -93
rect 357 -94 358 -93
rect 358 -94 359 -93
rect 359 -94 360 -93
rect 360 -94 361 -93
rect 361 -94 362 -93
rect 362 -94 363 -93
rect 363 -94 364 -93
rect 364 -94 365 -93
rect 365 -94 366 -93
rect 366 -94 367 -93
rect 367 -94 368 -93
rect 368 -94 369 -93
rect 369 -94 370 -93
rect 370 -94 371 -93
rect 371 -94 372 -93
rect 372 -94 373 -93
rect 373 -94 374 -93
rect 374 -94 375 -93
rect 375 -94 376 -93
rect 376 -94 377 -93
rect 377 -94 378 -93
rect 378 -94 379 -93
rect 379 -94 380 -93
rect 380 -94 381 -93
rect 381 -94 382 -93
rect 382 -94 383 -93
rect 383 -94 384 -93
rect 384 -94 385 -93
rect 385 -94 386 -93
rect 386 -94 387 -93
rect 387 -94 388 -93
rect 388 -94 389 -93
rect 389 -94 390 -93
rect 390 -94 391 -93
rect 391 -94 392 -93
rect 392 -94 393 -93
rect 393 -94 394 -93
rect 394 -94 395 -93
rect 395 -94 396 -93
rect 396 -94 397 -93
rect 397 -94 398 -93
rect 398 -94 399 -93
rect 399 -94 400 -93
rect 400 -94 401 -93
rect 401 -94 402 -93
rect 402 -94 403 -93
rect 403 -94 404 -93
rect 404 -94 405 -93
rect 405 -94 406 -93
rect 406 -94 407 -93
rect 407 -94 408 -93
rect 408 -94 409 -93
rect 409 -94 410 -93
rect 410 -94 411 -93
rect 411 -94 412 -93
rect 412 -94 413 -93
rect 413 -94 414 -93
rect 414 -94 415 -93
rect 415 -94 416 -93
rect 416 -94 417 -93
rect 417 -94 418 -93
rect 418 -94 419 -93
rect 419 -94 420 -93
rect 420 -94 421 -93
rect 421 -94 422 -93
rect 422 -94 423 -93
rect 423 -94 424 -93
rect 424 -94 425 -93
rect 425 -94 426 -93
rect 426 -94 427 -93
rect 427 -94 428 -93
rect 428 -94 429 -93
rect 429 -94 430 -93
rect 430 -94 431 -93
rect 431 -94 432 -93
rect 432 -94 433 -93
rect 433 -94 434 -93
rect 434 -94 435 -93
rect 435 -94 436 -93
rect 436 -94 437 -93
rect 437 -94 438 -93
rect 438 -94 439 -93
rect 439 -94 440 -93
rect 440 -94 441 -93
rect 441 -94 442 -93
rect 442 -94 443 -93
rect 443 -94 444 -93
rect 444 -94 445 -93
rect 445 -94 446 -93
rect 446 -94 447 -93
rect 447 -94 448 -93
rect 448 -94 449 -93
rect 449 -94 450 -93
rect 450 -94 451 -93
rect 451 -94 452 -93
rect 452 -94 453 -93
rect 453 -94 454 -93
rect 454 -94 455 -93
rect 455 -94 456 -93
rect 456 -94 457 -93
rect 457 -94 458 -93
rect 458 -94 459 -93
rect 459 -94 460 -93
rect 460 -94 461 -93
rect 461 -94 462 -93
rect 462 -94 463 -93
rect 463 -94 464 -93
rect 464 -94 465 -93
rect 465 -94 466 -93
rect 466 -94 467 -93
rect 467 -94 468 -93
rect 468 -94 469 -93
rect 469 -94 470 -93
rect 470 -94 471 -93
rect 471 -94 472 -93
rect 472 -94 473 -93
rect 473 -94 474 -93
rect 474 -94 475 -93
rect 475 -94 476 -93
rect 476 -94 477 -93
rect 477 -94 478 -93
rect 478 -94 479 -93
rect 479 -94 480 -93
rect 2 -95 3 -94
rect 3 -95 4 -94
rect 4 -95 5 -94
rect 5 -95 6 -94
rect 6 -95 7 -94
rect 7 -95 8 -94
rect 8 -95 9 -94
rect 9 -95 10 -94
rect 10 -95 11 -94
rect 23 -95 24 -94
rect 24 -95 25 -94
rect 25 -95 26 -94
rect 26 -95 27 -94
rect 27 -95 28 -94
rect 28 -95 29 -94
rect 29 -95 30 -94
rect 30 -95 31 -94
rect 31 -95 32 -94
rect 32 -95 33 -94
rect 33 -95 34 -94
rect 34 -95 35 -94
rect 35 -95 36 -94
rect 36 -95 37 -94
rect 37 -95 38 -94
rect 38 -95 39 -94
rect 39 -95 40 -94
rect 40 -95 41 -94
rect 41 -95 42 -94
rect 42 -95 43 -94
rect 55 -95 56 -94
rect 56 -95 57 -94
rect 57 -95 58 -94
rect 58 -95 59 -94
rect 59 -95 60 -94
rect 60 -95 61 -94
rect 61 -95 62 -94
rect 62 -95 63 -94
rect 63 -95 64 -94
rect 64 -95 65 -94
rect 65 -95 66 -94
rect 66 -95 67 -94
rect 67 -95 68 -94
rect 68 -95 69 -94
rect 69 -95 70 -94
rect 70 -95 71 -94
rect 71 -95 72 -94
rect 72 -95 73 -94
rect 73 -95 74 -94
rect 74 -95 75 -94
rect 87 -95 88 -94
rect 88 -95 89 -94
rect 89 -95 90 -94
rect 90 -95 91 -94
rect 91 -95 92 -94
rect 92 -95 93 -94
rect 93 -95 94 -94
rect 94 -95 95 -94
rect 95 -95 96 -94
rect 96 -95 97 -94
rect 97 -95 98 -94
rect 98 -95 99 -94
rect 99 -95 100 -94
rect 100 -95 101 -94
rect 101 -95 102 -94
rect 102 -95 103 -94
rect 103 -95 104 -94
rect 104 -95 105 -94
rect 105 -95 106 -94
rect 106 -95 107 -94
rect 119 -95 120 -94
rect 120 -95 121 -94
rect 121 -95 122 -94
rect 122 -95 123 -94
rect 123 -95 124 -94
rect 124 -95 125 -94
rect 125 -95 126 -94
rect 126 -95 127 -94
rect 127 -95 128 -94
rect 128 -95 129 -94
rect 129 -95 130 -94
rect 130 -95 131 -94
rect 131 -95 132 -94
rect 132 -95 133 -94
rect 133 -95 134 -94
rect 134 -95 135 -94
rect 135 -95 136 -94
rect 136 -95 137 -94
rect 137 -95 138 -94
rect 138 -95 139 -94
rect 151 -95 152 -94
rect 152 -95 153 -94
rect 153 -95 154 -94
rect 154 -95 155 -94
rect 155 -95 156 -94
rect 156 -95 157 -94
rect 157 -95 158 -94
rect 158 -95 159 -94
rect 159 -95 160 -94
rect 160 -95 161 -94
rect 161 -95 162 -94
rect 162 -95 163 -94
rect 163 -95 164 -94
rect 164 -95 165 -94
rect 165 -95 166 -94
rect 166 -95 167 -94
rect 167 -95 168 -94
rect 168 -95 169 -94
rect 169 -95 170 -94
rect 170 -95 171 -94
rect 183 -95 184 -94
rect 184 -95 185 -94
rect 185 -95 186 -94
rect 186 -95 187 -94
rect 187 -95 188 -94
rect 188 -95 189 -94
rect 189 -95 190 -94
rect 190 -95 191 -94
rect 191 -95 192 -94
rect 192 -95 193 -94
rect 193 -95 194 -94
rect 194 -95 195 -94
rect 195 -95 196 -94
rect 196 -95 197 -94
rect 197 -95 198 -94
rect 198 -95 199 -94
rect 199 -95 200 -94
rect 200 -95 201 -94
rect 201 -95 202 -94
rect 202 -95 203 -94
rect 203 -95 204 -94
rect 204 -95 205 -94
rect 205 -95 206 -94
rect 206 -95 207 -94
rect 207 -95 208 -94
rect 208 -95 209 -94
rect 209 -95 210 -94
rect 210 -95 211 -94
rect 211 -95 212 -94
rect 212 -95 213 -94
rect 213 -95 214 -94
rect 214 -95 215 -94
rect 215 -95 216 -94
rect 216 -95 217 -94
rect 217 -95 218 -94
rect 218 -95 219 -94
rect 219 -95 220 -94
rect 220 -95 221 -94
rect 221 -95 222 -94
rect 222 -95 223 -94
rect 223 -95 224 -94
rect 224 -95 225 -94
rect 225 -95 226 -94
rect 226 -95 227 -94
rect 227 -95 228 -94
rect 228 -95 229 -94
rect 229 -95 230 -94
rect 230 -95 231 -94
rect 231 -95 232 -94
rect 232 -95 233 -94
rect 233 -95 234 -94
rect 234 -95 235 -94
rect 235 -95 236 -94
rect 236 -95 237 -94
rect 237 -95 238 -94
rect 238 -95 239 -94
rect 239 -95 240 -94
rect 240 -95 241 -94
rect 241 -95 242 -94
rect 242 -95 243 -94
rect 243 -95 244 -94
rect 244 -95 245 -94
rect 245 -95 246 -94
rect 246 -95 247 -94
rect 247 -95 248 -94
rect 248 -95 249 -94
rect 249 -95 250 -94
rect 250 -95 251 -94
rect 251 -95 252 -94
rect 252 -95 253 -94
rect 253 -95 254 -94
rect 254 -95 255 -94
rect 255 -95 256 -94
rect 256 -95 257 -94
rect 257 -95 258 -94
rect 258 -95 259 -94
rect 259 -95 260 -94
rect 260 -95 261 -94
rect 261 -95 262 -94
rect 262 -95 263 -94
rect 263 -95 264 -94
rect 264 -95 265 -94
rect 265 -95 266 -94
rect 266 -95 267 -94
rect 267 -95 268 -94
rect 268 -95 269 -94
rect 269 -95 270 -94
rect 270 -95 271 -94
rect 271 -95 272 -94
rect 272 -95 273 -94
rect 273 -95 274 -94
rect 274 -95 275 -94
rect 275 -95 276 -94
rect 276 -95 277 -94
rect 277 -95 278 -94
rect 278 -95 279 -94
rect 279 -95 280 -94
rect 280 -95 281 -94
rect 281 -95 282 -94
rect 282 -95 283 -94
rect 283 -95 284 -94
rect 284 -95 285 -94
rect 285 -95 286 -94
rect 286 -95 287 -94
rect 287 -95 288 -94
rect 288 -95 289 -94
rect 289 -95 290 -94
rect 290 -95 291 -94
rect 291 -95 292 -94
rect 292 -95 293 -94
rect 293 -95 294 -94
rect 294 -95 295 -94
rect 295 -95 296 -94
rect 296 -95 297 -94
rect 297 -95 298 -94
rect 298 -95 299 -94
rect 299 -95 300 -94
rect 300 -95 301 -94
rect 301 -95 302 -94
rect 302 -95 303 -94
rect 303 -95 304 -94
rect 304 -95 305 -94
rect 305 -95 306 -94
rect 306 -95 307 -94
rect 307 -95 308 -94
rect 308 -95 309 -94
rect 309 -95 310 -94
rect 310 -95 311 -94
rect 311 -95 312 -94
rect 312 -95 313 -94
rect 313 -95 314 -94
rect 314 -95 315 -94
rect 315 -95 316 -94
rect 316 -95 317 -94
rect 317 -95 318 -94
rect 318 -95 319 -94
rect 319 -95 320 -94
rect 320 -95 321 -94
rect 321 -95 322 -94
rect 322 -95 323 -94
rect 323 -95 324 -94
rect 324 -95 325 -94
rect 325 -95 326 -94
rect 326 -95 327 -94
rect 327 -95 328 -94
rect 328 -95 329 -94
rect 329 -95 330 -94
rect 330 -95 331 -94
rect 331 -95 332 -94
rect 332 -95 333 -94
rect 333 -95 334 -94
rect 334 -95 335 -94
rect 335 -95 336 -94
rect 336 -95 337 -94
rect 337 -95 338 -94
rect 338 -95 339 -94
rect 339 -95 340 -94
rect 340 -95 341 -94
rect 341 -95 342 -94
rect 342 -95 343 -94
rect 343 -95 344 -94
rect 344 -95 345 -94
rect 345 -95 346 -94
rect 346 -95 347 -94
rect 347 -95 348 -94
rect 348 -95 349 -94
rect 349 -95 350 -94
rect 350 -95 351 -94
rect 351 -95 352 -94
rect 352 -95 353 -94
rect 353 -95 354 -94
rect 354 -95 355 -94
rect 355 -95 356 -94
rect 356 -95 357 -94
rect 357 -95 358 -94
rect 358 -95 359 -94
rect 359 -95 360 -94
rect 360 -95 361 -94
rect 361 -95 362 -94
rect 362 -95 363 -94
rect 363 -95 364 -94
rect 364 -95 365 -94
rect 365 -95 366 -94
rect 366 -95 367 -94
rect 367 -95 368 -94
rect 368 -95 369 -94
rect 369 -95 370 -94
rect 370 -95 371 -94
rect 371 -95 372 -94
rect 372 -95 373 -94
rect 373 -95 374 -94
rect 374 -95 375 -94
rect 375 -95 376 -94
rect 376 -95 377 -94
rect 377 -95 378 -94
rect 378 -95 379 -94
rect 379 -95 380 -94
rect 380 -95 381 -94
rect 381 -95 382 -94
rect 382 -95 383 -94
rect 383 -95 384 -94
rect 384 -95 385 -94
rect 385 -95 386 -94
rect 386 -95 387 -94
rect 387 -95 388 -94
rect 388 -95 389 -94
rect 389 -95 390 -94
rect 390 -95 391 -94
rect 391 -95 392 -94
rect 392 -95 393 -94
rect 393 -95 394 -94
rect 394 -95 395 -94
rect 395 -95 396 -94
rect 396 -95 397 -94
rect 397 -95 398 -94
rect 398 -95 399 -94
rect 399 -95 400 -94
rect 400 -95 401 -94
rect 401 -95 402 -94
rect 402 -95 403 -94
rect 403 -95 404 -94
rect 404 -95 405 -94
rect 405 -95 406 -94
rect 406 -95 407 -94
rect 407 -95 408 -94
rect 408 -95 409 -94
rect 409 -95 410 -94
rect 410 -95 411 -94
rect 411 -95 412 -94
rect 412 -95 413 -94
rect 413 -95 414 -94
rect 414 -95 415 -94
rect 415 -95 416 -94
rect 416 -95 417 -94
rect 417 -95 418 -94
rect 418 -95 419 -94
rect 419 -95 420 -94
rect 420 -95 421 -94
rect 421 -95 422 -94
rect 422 -95 423 -94
rect 423 -95 424 -94
rect 424 -95 425 -94
rect 425 -95 426 -94
rect 426 -95 427 -94
rect 427 -95 428 -94
rect 428 -95 429 -94
rect 429 -95 430 -94
rect 430 -95 431 -94
rect 431 -95 432 -94
rect 432 -95 433 -94
rect 433 -95 434 -94
rect 434 -95 435 -94
rect 435 -95 436 -94
rect 436 -95 437 -94
rect 437 -95 438 -94
rect 438 -95 439 -94
rect 439 -95 440 -94
rect 440 -95 441 -94
rect 441 -95 442 -94
rect 442 -95 443 -94
rect 443 -95 444 -94
rect 444 -95 445 -94
rect 445 -95 446 -94
rect 446 -95 447 -94
rect 447 -95 448 -94
rect 448 -95 449 -94
rect 449 -95 450 -94
rect 450 -95 451 -94
rect 451 -95 452 -94
rect 452 -95 453 -94
rect 453 -95 454 -94
rect 454 -95 455 -94
rect 455 -95 456 -94
rect 456 -95 457 -94
rect 457 -95 458 -94
rect 458 -95 459 -94
rect 459 -95 460 -94
rect 460 -95 461 -94
rect 461 -95 462 -94
rect 462 -95 463 -94
rect 463 -95 464 -94
rect 464 -95 465 -94
rect 465 -95 466 -94
rect 466 -95 467 -94
rect 467 -95 468 -94
rect 468 -95 469 -94
rect 469 -95 470 -94
rect 470 -95 471 -94
rect 471 -95 472 -94
rect 472 -95 473 -94
rect 473 -95 474 -94
rect 474 -95 475 -94
rect 475 -95 476 -94
rect 476 -95 477 -94
rect 477 -95 478 -94
rect 478 -95 479 -94
rect 479 -95 480 -94
rect 2 -96 3 -95
rect 3 -96 4 -95
rect 4 -96 5 -95
rect 5 -96 6 -95
rect 6 -96 7 -95
rect 7 -96 8 -95
rect 8 -96 9 -95
rect 9 -96 10 -95
rect 10 -96 11 -95
rect 11 -96 12 -95
rect 21 -96 22 -95
rect 22 -96 23 -95
rect 23 -96 24 -95
rect 24 -96 25 -95
rect 25 -96 26 -95
rect 26 -96 27 -95
rect 27 -96 28 -95
rect 28 -96 29 -95
rect 29 -96 30 -95
rect 30 -96 31 -95
rect 31 -96 32 -95
rect 32 -96 33 -95
rect 33 -96 34 -95
rect 34 -96 35 -95
rect 35 -96 36 -95
rect 36 -96 37 -95
rect 37 -96 38 -95
rect 38 -96 39 -95
rect 39 -96 40 -95
rect 40 -96 41 -95
rect 41 -96 42 -95
rect 42 -96 43 -95
rect 43 -96 44 -95
rect 54 -96 55 -95
rect 55 -96 56 -95
rect 56 -96 57 -95
rect 57 -96 58 -95
rect 58 -96 59 -95
rect 59 -96 60 -95
rect 60 -96 61 -95
rect 61 -96 62 -95
rect 62 -96 63 -95
rect 63 -96 64 -95
rect 64 -96 65 -95
rect 65 -96 66 -95
rect 66 -96 67 -95
rect 67 -96 68 -95
rect 68 -96 69 -95
rect 69 -96 70 -95
rect 70 -96 71 -95
rect 71 -96 72 -95
rect 72 -96 73 -95
rect 73 -96 74 -95
rect 74 -96 75 -95
rect 75 -96 76 -95
rect 85 -96 86 -95
rect 86 -96 87 -95
rect 87 -96 88 -95
rect 88 -96 89 -95
rect 89 -96 90 -95
rect 90 -96 91 -95
rect 91 -96 92 -95
rect 92 -96 93 -95
rect 93 -96 94 -95
rect 94 -96 95 -95
rect 95 -96 96 -95
rect 96 -96 97 -95
rect 97 -96 98 -95
rect 98 -96 99 -95
rect 99 -96 100 -95
rect 100 -96 101 -95
rect 101 -96 102 -95
rect 102 -96 103 -95
rect 103 -96 104 -95
rect 104 -96 105 -95
rect 105 -96 106 -95
rect 106 -96 107 -95
rect 107 -96 108 -95
rect 118 -96 119 -95
rect 119 -96 120 -95
rect 120 -96 121 -95
rect 121 -96 122 -95
rect 122 -96 123 -95
rect 123 -96 124 -95
rect 124 -96 125 -95
rect 125 -96 126 -95
rect 126 -96 127 -95
rect 127 -96 128 -95
rect 128 -96 129 -95
rect 129 -96 130 -95
rect 130 -96 131 -95
rect 131 -96 132 -95
rect 132 -96 133 -95
rect 133 -96 134 -95
rect 134 -96 135 -95
rect 135 -96 136 -95
rect 136 -96 137 -95
rect 137 -96 138 -95
rect 138 -96 139 -95
rect 139 -96 140 -95
rect 149 -96 150 -95
rect 150 -96 151 -95
rect 151 -96 152 -95
rect 152 -96 153 -95
rect 153 -96 154 -95
rect 154 -96 155 -95
rect 155 -96 156 -95
rect 156 -96 157 -95
rect 157 -96 158 -95
rect 158 -96 159 -95
rect 159 -96 160 -95
rect 160 -96 161 -95
rect 161 -96 162 -95
rect 162 -96 163 -95
rect 163 -96 164 -95
rect 164 -96 165 -95
rect 165 -96 166 -95
rect 166 -96 167 -95
rect 167 -96 168 -95
rect 168 -96 169 -95
rect 169 -96 170 -95
rect 170 -96 171 -95
rect 171 -96 172 -95
rect 181 -96 182 -95
rect 182 -96 183 -95
rect 183 -96 184 -95
rect 184 -96 185 -95
rect 185 -96 186 -95
rect 186 -96 187 -95
rect 187 -96 188 -95
rect 188 -96 189 -95
rect 189 -96 190 -95
rect 190 -96 191 -95
rect 191 -96 192 -95
rect 2 -97 3 -96
rect 3 -97 4 -96
rect 4 -97 5 -96
rect 5 -97 6 -96
rect 6 -97 7 -96
rect 7 -97 8 -96
rect 8 -97 9 -96
rect 9 -97 10 -96
rect 10 -97 11 -96
rect 11 -97 12 -96
rect 21 -97 22 -96
rect 22 -97 23 -96
rect 23 -97 24 -96
rect 24 -97 25 -96
rect 25 -97 26 -96
rect 26 -97 27 -96
rect 27 -97 28 -96
rect 28 -97 29 -96
rect 29 -97 30 -96
rect 30 -97 31 -96
rect 31 -97 32 -96
rect 32 -97 33 -96
rect 33 -97 34 -96
rect 34 -97 35 -96
rect 35 -97 36 -96
rect 36 -97 37 -96
rect 37 -97 38 -96
rect 38 -97 39 -96
rect 39 -97 40 -96
rect 40 -97 41 -96
rect 41 -97 42 -96
rect 42 -97 43 -96
rect 43 -97 44 -96
rect 53 -97 54 -96
rect 54 -97 55 -96
rect 55 -97 56 -96
rect 56 -97 57 -96
rect 57 -97 58 -96
rect 58 -97 59 -96
rect 59 -97 60 -96
rect 60 -97 61 -96
rect 61 -97 62 -96
rect 62 -97 63 -96
rect 63 -97 64 -96
rect 64 -97 65 -96
rect 65 -97 66 -96
rect 66 -97 67 -96
rect 67 -97 68 -96
rect 68 -97 69 -96
rect 69 -97 70 -96
rect 70 -97 71 -96
rect 71 -97 72 -96
rect 72 -97 73 -96
rect 73 -97 74 -96
rect 74 -97 75 -96
rect 75 -97 76 -96
rect 85 -97 86 -96
rect 86 -97 87 -96
rect 87 -97 88 -96
rect 88 -97 89 -96
rect 89 -97 90 -96
rect 90 -97 91 -96
rect 91 -97 92 -96
rect 92 -97 93 -96
rect 93 -97 94 -96
rect 94 -97 95 -96
rect 95 -97 96 -96
rect 96 -97 97 -96
rect 97 -97 98 -96
rect 98 -97 99 -96
rect 99 -97 100 -96
rect 100 -97 101 -96
rect 101 -97 102 -96
rect 102 -97 103 -96
rect 103 -97 104 -96
rect 104 -97 105 -96
rect 105 -97 106 -96
rect 106 -97 107 -96
rect 107 -97 108 -96
rect 117 -97 118 -96
rect 118 -97 119 -96
rect 119 -97 120 -96
rect 120 -97 121 -96
rect 121 -97 122 -96
rect 122 -97 123 -96
rect 123 -97 124 -96
rect 124 -97 125 -96
rect 125 -97 126 -96
rect 126 -97 127 -96
rect 127 -97 128 -96
rect 128 -97 129 -96
rect 129 -97 130 -96
rect 130 -97 131 -96
rect 131 -97 132 -96
rect 132 -97 133 -96
rect 133 -97 134 -96
rect 134 -97 135 -96
rect 135 -97 136 -96
rect 136 -97 137 -96
rect 137 -97 138 -96
rect 138 -97 139 -96
rect 139 -97 140 -96
rect 149 -97 150 -96
rect 150 -97 151 -96
rect 151 -97 152 -96
rect 152 -97 153 -96
rect 153 -97 154 -96
rect 154 -97 155 -96
rect 155 -97 156 -96
rect 156 -97 157 -96
rect 157 -97 158 -96
rect 158 -97 159 -96
rect 159 -97 160 -96
rect 160 -97 161 -96
rect 161 -97 162 -96
rect 162 -97 163 -96
rect 163 -97 164 -96
rect 164 -97 165 -96
rect 165 -97 166 -96
rect 166 -97 167 -96
rect 167 -97 168 -96
rect 168 -97 169 -96
rect 169 -97 170 -96
rect 170 -97 171 -96
rect 171 -97 172 -96
rect 181 -97 182 -96
rect 182 -97 183 -96
rect 183 -97 184 -96
rect 184 -97 185 -96
rect 185 -97 186 -96
rect 186 -97 187 -96
rect 187 -97 188 -96
rect 188 -97 189 -96
rect 189 -97 190 -96
rect 190 -97 191 -96
rect 191 -97 192 -96
rect 2 -98 3 -97
rect 3 -98 4 -97
rect 4 -98 5 -97
rect 5 -98 6 -97
rect 6 -98 7 -97
rect 7 -98 8 -97
rect 8 -98 9 -97
rect 9 -98 10 -97
rect 10 -98 11 -97
rect 11 -98 12 -97
rect 21 -98 22 -97
rect 22 -98 23 -97
rect 23 -98 24 -97
rect 24 -98 25 -97
rect 25 -98 26 -97
rect 26 -98 27 -97
rect 27 -98 28 -97
rect 28 -98 29 -97
rect 29 -98 30 -97
rect 30 -98 31 -97
rect 31 -98 32 -97
rect 32 -98 33 -97
rect 33 -98 34 -97
rect 34 -98 35 -97
rect 35 -98 36 -97
rect 36 -98 37 -97
rect 37 -98 38 -97
rect 38 -98 39 -97
rect 39 -98 40 -97
rect 40 -98 41 -97
rect 41 -98 42 -97
rect 42 -98 43 -97
rect 43 -98 44 -97
rect 53 -98 54 -97
rect 54 -98 55 -97
rect 55 -98 56 -97
rect 56 -98 57 -97
rect 57 -98 58 -97
rect 58 -98 59 -97
rect 59 -98 60 -97
rect 60 -98 61 -97
rect 61 -98 62 -97
rect 62 -98 63 -97
rect 63 -98 64 -97
rect 64 -98 65 -97
rect 65 -98 66 -97
rect 66 -98 67 -97
rect 67 -98 68 -97
rect 68 -98 69 -97
rect 69 -98 70 -97
rect 70 -98 71 -97
rect 71 -98 72 -97
rect 72 -98 73 -97
rect 73 -98 74 -97
rect 74 -98 75 -97
rect 75 -98 76 -97
rect 85 -98 86 -97
rect 86 -98 87 -97
rect 87 -98 88 -97
rect 88 -98 89 -97
rect 89 -98 90 -97
rect 90 -98 91 -97
rect 91 -98 92 -97
rect 92 -98 93 -97
rect 93 -98 94 -97
rect 94 -98 95 -97
rect 95 -98 96 -97
rect 96 -98 97 -97
rect 97 -98 98 -97
rect 98 -98 99 -97
rect 99 -98 100 -97
rect 100 -98 101 -97
rect 101 -98 102 -97
rect 102 -98 103 -97
rect 103 -98 104 -97
rect 104 -98 105 -97
rect 105 -98 106 -97
rect 106 -98 107 -97
rect 107 -98 108 -97
rect 117 -98 118 -97
rect 118 -98 119 -97
rect 119 -98 120 -97
rect 120 -98 121 -97
rect 121 -98 122 -97
rect 122 -98 123 -97
rect 123 -98 124 -97
rect 124 -98 125 -97
rect 125 -98 126 -97
rect 126 -98 127 -97
rect 127 -98 128 -97
rect 128 -98 129 -97
rect 129 -98 130 -97
rect 130 -98 131 -97
rect 131 -98 132 -97
rect 132 -98 133 -97
rect 133 -98 134 -97
rect 134 -98 135 -97
rect 135 -98 136 -97
rect 136 -98 137 -97
rect 137 -98 138 -97
rect 138 -98 139 -97
rect 139 -98 140 -97
rect 149 -98 150 -97
rect 150 -98 151 -97
rect 151 -98 152 -97
rect 152 -98 153 -97
rect 153 -98 154 -97
rect 154 -98 155 -97
rect 155 -98 156 -97
rect 156 -98 157 -97
rect 157 -98 158 -97
rect 158 -98 159 -97
rect 159 -98 160 -97
rect 160 -98 161 -97
rect 161 -98 162 -97
rect 162 -98 163 -97
rect 163 -98 164 -97
rect 164 -98 165 -97
rect 165 -98 166 -97
rect 166 -98 167 -97
rect 167 -98 168 -97
rect 168 -98 169 -97
rect 169 -98 170 -97
rect 170 -98 171 -97
rect 171 -98 172 -97
rect 181 -98 182 -97
rect 182 -98 183 -97
rect 183 -98 184 -97
rect 184 -98 185 -97
rect 185 -98 186 -97
rect 186 -98 187 -97
rect 187 -98 188 -97
rect 188 -98 189 -97
rect 189 -98 190 -97
rect 190 -98 191 -97
rect 191 -98 192 -97
rect 2 -99 3 -98
rect 3 -99 4 -98
rect 4 -99 5 -98
rect 5 -99 6 -98
rect 6 -99 7 -98
rect 7 -99 8 -98
rect 8 -99 9 -98
rect 9 -99 10 -98
rect 10 -99 11 -98
rect 11 -99 12 -98
rect 22 -99 23 -98
rect 23 -99 24 -98
rect 24 -99 25 -98
rect 25 -99 26 -98
rect 26 -99 27 -98
rect 27 -99 28 -98
rect 28 -99 29 -98
rect 29 -99 30 -98
rect 30 -99 31 -98
rect 31 -99 32 -98
rect 32 -99 33 -98
rect 33 -99 34 -98
rect 34 -99 35 -98
rect 35 -99 36 -98
rect 36 -99 37 -98
rect 37 -99 38 -98
rect 38 -99 39 -98
rect 39 -99 40 -98
rect 40 -99 41 -98
rect 41 -99 42 -98
rect 42 -99 43 -98
rect 43 -99 44 -98
rect 54 -99 55 -98
rect 55 -99 56 -98
rect 56 -99 57 -98
rect 57 -99 58 -98
rect 58 -99 59 -98
rect 59 -99 60 -98
rect 60 -99 61 -98
rect 61 -99 62 -98
rect 62 -99 63 -98
rect 63 -99 64 -98
rect 64 -99 65 -98
rect 65 -99 66 -98
rect 66 -99 67 -98
rect 67 -99 68 -98
rect 68 -99 69 -98
rect 69 -99 70 -98
rect 70 -99 71 -98
rect 71 -99 72 -98
rect 72 -99 73 -98
rect 73 -99 74 -98
rect 74 -99 75 -98
rect 75 -99 76 -98
rect 86 -99 87 -98
rect 87 -99 88 -98
rect 88 -99 89 -98
rect 89 -99 90 -98
rect 90 -99 91 -98
rect 91 -99 92 -98
rect 92 -99 93 -98
rect 93 -99 94 -98
rect 94 -99 95 -98
rect 95 -99 96 -98
rect 96 -99 97 -98
rect 97 -99 98 -98
rect 98 -99 99 -98
rect 99 -99 100 -98
rect 100 -99 101 -98
rect 101 -99 102 -98
rect 102 -99 103 -98
rect 103 -99 104 -98
rect 104 -99 105 -98
rect 105 -99 106 -98
rect 106 -99 107 -98
rect 107 -99 108 -98
rect 118 -99 119 -98
rect 119 -99 120 -98
rect 120 -99 121 -98
rect 121 -99 122 -98
rect 122 -99 123 -98
rect 123 -99 124 -98
rect 124 -99 125 -98
rect 125 -99 126 -98
rect 126 -99 127 -98
rect 127 -99 128 -98
rect 128 -99 129 -98
rect 129 -99 130 -98
rect 130 -99 131 -98
rect 131 -99 132 -98
rect 132 -99 133 -98
rect 133 -99 134 -98
rect 134 -99 135 -98
rect 135 -99 136 -98
rect 136 -99 137 -98
rect 137 -99 138 -98
rect 138 -99 139 -98
rect 139 -99 140 -98
rect 150 -99 151 -98
rect 151 -99 152 -98
rect 152 -99 153 -98
rect 153 -99 154 -98
rect 154 -99 155 -98
rect 155 -99 156 -98
rect 156 -99 157 -98
rect 157 -99 158 -98
rect 158 -99 159 -98
rect 159 -99 160 -98
rect 160 -99 161 -98
rect 161 -99 162 -98
rect 162 -99 163 -98
rect 163 -99 164 -98
rect 164 -99 165 -98
rect 165 -99 166 -98
rect 166 -99 167 -98
rect 167 -99 168 -98
rect 168 -99 169 -98
rect 169 -99 170 -98
rect 170 -99 171 -98
rect 171 -99 172 -98
rect 182 -99 183 -98
rect 183 -99 184 -98
rect 184 -99 185 -98
rect 185 -99 186 -98
rect 186 -99 187 -98
rect 187 -99 188 -98
rect 188 -99 189 -98
rect 189 -99 190 -98
rect 190 -99 191 -98
rect 191 -99 192 -98
rect 2 -100 3 -99
rect 3 -100 4 -99
rect 4 -100 5 -99
rect 5 -100 6 -99
rect 6 -100 7 -99
rect 7 -100 8 -99
rect 8 -100 9 -99
rect 9 -100 10 -99
rect 10 -100 11 -99
rect 11 -100 12 -99
rect 16 -100 17 -99
rect 17 -100 18 -99
rect 22 -100 23 -99
rect 23 -100 24 -99
rect 24 -100 25 -99
rect 25 -100 26 -99
rect 26 -100 27 -99
rect 27 -100 28 -99
rect 28 -100 29 -99
rect 29 -100 30 -99
rect 30 -100 31 -99
rect 31 -100 32 -99
rect 32 -100 33 -99
rect 33 -100 34 -99
rect 34 -100 35 -99
rect 35 -100 36 -99
rect 36 -100 37 -99
rect 37 -100 38 -99
rect 38 -100 39 -99
rect 39 -100 40 -99
rect 40 -100 41 -99
rect 41 -100 42 -99
rect 42 -100 43 -99
rect 43 -100 44 -99
rect 48 -100 49 -99
rect 49 -100 50 -99
rect 54 -100 55 -99
rect 55 -100 56 -99
rect 56 -100 57 -99
rect 57 -100 58 -99
rect 58 -100 59 -99
rect 59 -100 60 -99
rect 60 -100 61 -99
rect 61 -100 62 -99
rect 62 -100 63 -99
rect 63 -100 64 -99
rect 64 -100 65 -99
rect 65 -100 66 -99
rect 66 -100 67 -99
rect 67 -100 68 -99
rect 68 -100 69 -99
rect 69 -100 70 -99
rect 70 -100 71 -99
rect 71 -100 72 -99
rect 72 -100 73 -99
rect 73 -100 74 -99
rect 74 -100 75 -99
rect 75 -100 76 -99
rect 80 -100 81 -99
rect 81 -100 82 -99
rect 86 -100 87 -99
rect 87 -100 88 -99
rect 88 -100 89 -99
rect 89 -100 90 -99
rect 90 -100 91 -99
rect 91 -100 92 -99
rect 92 -100 93 -99
rect 93 -100 94 -99
rect 94 -100 95 -99
rect 95 -100 96 -99
rect 96 -100 97 -99
rect 97 -100 98 -99
rect 98 -100 99 -99
rect 99 -100 100 -99
rect 100 -100 101 -99
rect 101 -100 102 -99
rect 102 -100 103 -99
rect 103 -100 104 -99
rect 104 -100 105 -99
rect 105 -100 106 -99
rect 106 -100 107 -99
rect 107 -100 108 -99
rect 112 -100 113 -99
rect 113 -100 114 -99
rect 118 -100 119 -99
rect 119 -100 120 -99
rect 120 -100 121 -99
rect 121 -100 122 -99
rect 122 -100 123 -99
rect 123 -100 124 -99
rect 124 -100 125 -99
rect 125 -100 126 -99
rect 126 -100 127 -99
rect 127 -100 128 -99
rect 128 -100 129 -99
rect 129 -100 130 -99
rect 130 -100 131 -99
rect 131 -100 132 -99
rect 132 -100 133 -99
rect 133 -100 134 -99
rect 134 -100 135 -99
rect 135 -100 136 -99
rect 136 -100 137 -99
rect 137 -100 138 -99
rect 138 -100 139 -99
rect 139 -100 140 -99
rect 144 -100 145 -99
rect 145 -100 146 -99
rect 150 -100 151 -99
rect 151 -100 152 -99
rect 152 -100 153 -99
rect 153 -100 154 -99
rect 154 -100 155 -99
rect 155 -100 156 -99
rect 156 -100 157 -99
rect 157 -100 158 -99
rect 158 -100 159 -99
rect 159 -100 160 -99
rect 160 -100 161 -99
rect 161 -100 162 -99
rect 162 -100 163 -99
rect 163 -100 164 -99
rect 164 -100 165 -99
rect 165 -100 166 -99
rect 166 -100 167 -99
rect 167 -100 168 -99
rect 168 -100 169 -99
rect 169 -100 170 -99
rect 170 -100 171 -99
rect 171 -100 172 -99
rect 176 -100 177 -99
rect 177 -100 178 -99
rect 182 -100 183 -99
rect 183 -100 184 -99
rect 184 -100 185 -99
rect 185 -100 186 -99
rect 186 -100 187 -99
rect 187 -100 188 -99
rect 188 -100 189 -99
rect 189 -100 190 -99
rect 190 -100 191 -99
rect 191 -100 192 -99
rect 2 -101 3 -100
rect 3 -101 4 -100
rect 4 -101 5 -100
rect 5 -101 6 -100
rect 6 -101 7 -100
rect 7 -101 8 -100
rect 8 -101 9 -100
rect 9 -101 10 -100
rect 10 -101 11 -100
rect 11 -101 12 -100
rect 14 -101 15 -100
rect 15 -101 16 -100
rect 16 -101 17 -100
rect 17 -101 18 -100
rect 18 -101 19 -100
rect 22 -101 23 -100
rect 23 -101 24 -100
rect 24 -101 25 -100
rect 25 -101 26 -100
rect 26 -101 27 -100
rect 27 -101 28 -100
rect 28 -101 29 -100
rect 29 -101 30 -100
rect 30 -101 31 -100
rect 31 -101 32 -100
rect 34 -101 35 -100
rect 35 -101 36 -100
rect 36 -101 37 -100
rect 37 -101 38 -100
rect 38 -101 39 -100
rect 39 -101 40 -100
rect 40 -101 41 -100
rect 41 -101 42 -100
rect 42 -101 43 -100
rect 43 -101 44 -100
rect 46 -101 47 -100
rect 47 -101 48 -100
rect 48 -101 49 -100
rect 49 -101 50 -100
rect 50 -101 51 -100
rect 54 -101 55 -100
rect 55 -101 56 -100
rect 56 -101 57 -100
rect 57 -101 58 -100
rect 58 -101 59 -100
rect 59 -101 60 -100
rect 60 -101 61 -100
rect 61 -101 62 -100
rect 62 -101 63 -100
rect 63 -101 64 -100
rect 66 -101 67 -100
rect 67 -101 68 -100
rect 68 -101 69 -100
rect 69 -101 70 -100
rect 70 -101 71 -100
rect 71 -101 72 -100
rect 72 -101 73 -100
rect 73 -101 74 -100
rect 74 -101 75 -100
rect 75 -101 76 -100
rect 78 -101 79 -100
rect 79 -101 80 -100
rect 80 -101 81 -100
rect 81 -101 82 -100
rect 82 -101 83 -100
rect 86 -101 87 -100
rect 87 -101 88 -100
rect 88 -101 89 -100
rect 89 -101 90 -100
rect 90 -101 91 -100
rect 91 -101 92 -100
rect 92 -101 93 -100
rect 93 -101 94 -100
rect 94 -101 95 -100
rect 95 -101 96 -100
rect 98 -101 99 -100
rect 99 -101 100 -100
rect 100 -101 101 -100
rect 101 -101 102 -100
rect 102 -101 103 -100
rect 103 -101 104 -100
rect 104 -101 105 -100
rect 105 -101 106 -100
rect 106 -101 107 -100
rect 107 -101 108 -100
rect 110 -101 111 -100
rect 111 -101 112 -100
rect 112 -101 113 -100
rect 113 -101 114 -100
rect 114 -101 115 -100
rect 118 -101 119 -100
rect 119 -101 120 -100
rect 120 -101 121 -100
rect 121 -101 122 -100
rect 122 -101 123 -100
rect 123 -101 124 -100
rect 124 -101 125 -100
rect 125 -101 126 -100
rect 126 -101 127 -100
rect 127 -101 128 -100
rect 130 -101 131 -100
rect 131 -101 132 -100
rect 132 -101 133 -100
rect 133 -101 134 -100
rect 134 -101 135 -100
rect 135 -101 136 -100
rect 136 -101 137 -100
rect 137 -101 138 -100
rect 138 -101 139 -100
rect 139 -101 140 -100
rect 142 -101 143 -100
rect 143 -101 144 -100
rect 144 -101 145 -100
rect 145 -101 146 -100
rect 146 -101 147 -100
rect 150 -101 151 -100
rect 151 -101 152 -100
rect 152 -101 153 -100
rect 153 -101 154 -100
rect 154 -101 155 -100
rect 155 -101 156 -100
rect 156 -101 157 -100
rect 157 -101 158 -100
rect 158 -101 159 -100
rect 159 -101 160 -100
rect 162 -101 163 -100
rect 163 -101 164 -100
rect 164 -101 165 -100
rect 165 -101 166 -100
rect 166 -101 167 -100
rect 167 -101 168 -100
rect 168 -101 169 -100
rect 169 -101 170 -100
rect 170 -101 171 -100
rect 171 -101 172 -100
rect 174 -101 175 -100
rect 175 -101 176 -100
rect 176 -101 177 -100
rect 177 -101 178 -100
rect 178 -101 179 -100
rect 182 -101 183 -100
rect 183 -101 184 -100
rect 184 -101 185 -100
rect 185 -101 186 -100
rect 186 -101 187 -100
rect 187 -101 188 -100
rect 188 -101 189 -100
rect 189 -101 190 -100
rect 190 -101 191 -100
rect 191 -101 192 -100
rect 2 -102 3 -101
rect 3 -102 4 -101
rect 4 -102 5 -101
rect 5 -102 6 -101
rect 6 -102 7 -101
rect 7 -102 8 -101
rect 8 -102 9 -101
rect 9 -102 10 -101
rect 10 -102 11 -101
rect 11 -102 12 -101
rect 12 -102 13 -101
rect 13 -102 14 -101
rect 14 -102 15 -101
rect 15 -102 16 -101
rect 16 -102 17 -101
rect 17 -102 18 -101
rect 18 -102 19 -101
rect 19 -102 20 -101
rect 20 -102 21 -101
rect 21 -102 22 -101
rect 22 -102 23 -101
rect 23 -102 24 -101
rect 24 -102 25 -101
rect 25 -102 26 -101
rect 26 -102 27 -101
rect 27 -102 28 -101
rect 28 -102 29 -101
rect 29 -102 30 -101
rect 30 -102 31 -101
rect 34 -102 35 -101
rect 35 -102 36 -101
rect 36 -102 37 -101
rect 37 -102 38 -101
rect 38 -102 39 -101
rect 39 -102 40 -101
rect 40 -102 41 -101
rect 41 -102 42 -101
rect 42 -102 43 -101
rect 43 -102 44 -101
rect 44 -102 45 -101
rect 45 -102 46 -101
rect 46 -102 47 -101
rect 47 -102 48 -101
rect 48 -102 49 -101
rect 49 -102 50 -101
rect 50 -102 51 -101
rect 51 -102 52 -101
rect 52 -102 53 -101
rect 53 -102 54 -101
rect 54 -102 55 -101
rect 55 -102 56 -101
rect 56 -102 57 -101
rect 57 -102 58 -101
rect 58 -102 59 -101
rect 59 -102 60 -101
rect 60 -102 61 -101
rect 61 -102 62 -101
rect 62 -102 63 -101
rect 66 -102 67 -101
rect 67 -102 68 -101
rect 68 -102 69 -101
rect 69 -102 70 -101
rect 70 -102 71 -101
rect 71 -102 72 -101
rect 72 -102 73 -101
rect 73 -102 74 -101
rect 74 -102 75 -101
rect 75 -102 76 -101
rect 76 -102 77 -101
rect 77 -102 78 -101
rect 78 -102 79 -101
rect 79 -102 80 -101
rect 80 -102 81 -101
rect 81 -102 82 -101
rect 82 -102 83 -101
rect 83 -102 84 -101
rect 84 -102 85 -101
rect 85 -102 86 -101
rect 86 -102 87 -101
rect 87 -102 88 -101
rect 88 -102 89 -101
rect 89 -102 90 -101
rect 90 -102 91 -101
rect 91 -102 92 -101
rect 92 -102 93 -101
rect 93 -102 94 -101
rect 94 -102 95 -101
rect 98 -102 99 -101
rect 99 -102 100 -101
rect 100 -102 101 -101
rect 101 -102 102 -101
rect 102 -102 103 -101
rect 103 -102 104 -101
rect 104 -102 105 -101
rect 105 -102 106 -101
rect 106 -102 107 -101
rect 107 -102 108 -101
rect 108 -102 109 -101
rect 109 -102 110 -101
rect 110 -102 111 -101
rect 111 -102 112 -101
rect 112 -102 113 -101
rect 113 -102 114 -101
rect 114 -102 115 -101
rect 115 -102 116 -101
rect 116 -102 117 -101
rect 117 -102 118 -101
rect 118 -102 119 -101
rect 119 -102 120 -101
rect 120 -102 121 -101
rect 121 -102 122 -101
rect 122 -102 123 -101
rect 123 -102 124 -101
rect 124 -102 125 -101
rect 125 -102 126 -101
rect 126 -102 127 -101
rect 130 -102 131 -101
rect 131 -102 132 -101
rect 132 -102 133 -101
rect 133 -102 134 -101
rect 134 -102 135 -101
rect 135 -102 136 -101
rect 136 -102 137 -101
rect 137 -102 138 -101
rect 138 -102 139 -101
rect 139 -102 140 -101
rect 140 -102 141 -101
rect 141 -102 142 -101
rect 142 -102 143 -101
rect 143 -102 144 -101
rect 144 -102 145 -101
rect 145 -102 146 -101
rect 146 -102 147 -101
rect 147 -102 148 -101
rect 148 -102 149 -101
rect 149 -102 150 -101
rect 150 -102 151 -101
rect 151 -102 152 -101
rect 152 -102 153 -101
rect 153 -102 154 -101
rect 154 -102 155 -101
rect 155 -102 156 -101
rect 156 -102 157 -101
rect 157 -102 158 -101
rect 158 -102 159 -101
rect 162 -102 163 -101
rect 163 -102 164 -101
rect 164 -102 165 -101
rect 165 -102 166 -101
rect 166 -102 167 -101
rect 167 -102 168 -101
rect 168 -102 169 -101
rect 169 -102 170 -101
rect 170 -102 171 -101
rect 171 -102 172 -101
rect 172 -102 173 -101
rect 173 -102 174 -101
rect 174 -102 175 -101
rect 175 -102 176 -101
rect 176 -102 177 -101
rect 177 -102 178 -101
rect 178 -102 179 -101
rect 179 -102 180 -101
rect 180 -102 181 -101
rect 181 -102 182 -101
rect 182 -102 183 -101
rect 183 -102 184 -101
rect 184 -102 185 -101
rect 185 -102 186 -101
rect 186 -102 187 -101
rect 187 -102 188 -101
rect 188 -102 189 -101
rect 189 -102 190 -101
rect 190 -102 191 -101
rect 191 -102 192 -101
rect 2 -103 3 -102
rect 3 -103 4 -102
rect 4 -103 5 -102
rect 5 -103 6 -102
rect 6 -103 7 -102
rect 7 -103 8 -102
rect 8 -103 9 -102
rect 9 -103 10 -102
rect 10 -103 11 -102
rect 11 -103 12 -102
rect 12 -103 13 -102
rect 13 -103 14 -102
rect 14 -103 15 -102
rect 15 -103 16 -102
rect 16 -103 17 -102
rect 17 -103 18 -102
rect 18 -103 19 -102
rect 19 -103 20 -102
rect 20 -103 21 -102
rect 21 -103 22 -102
rect 22 -103 23 -102
rect 23 -103 24 -102
rect 24 -103 25 -102
rect 25 -103 26 -102
rect 26 -103 27 -102
rect 27 -103 28 -102
rect 28 -103 29 -102
rect 29 -103 30 -102
rect 30 -103 31 -102
rect 35 -103 36 -102
rect 36 -103 37 -102
rect 37 -103 38 -102
rect 38 -103 39 -102
rect 39 -103 40 -102
rect 40 -103 41 -102
rect 41 -103 42 -102
rect 42 -103 43 -102
rect 43 -103 44 -102
rect 44 -103 45 -102
rect 45 -103 46 -102
rect 46 -103 47 -102
rect 47 -103 48 -102
rect 48 -103 49 -102
rect 49 -103 50 -102
rect 50 -103 51 -102
rect 51 -103 52 -102
rect 52 -103 53 -102
rect 53 -103 54 -102
rect 54 -103 55 -102
rect 55 -103 56 -102
rect 56 -103 57 -102
rect 57 -103 58 -102
rect 58 -103 59 -102
rect 59 -103 60 -102
rect 60 -103 61 -102
rect 61 -103 62 -102
rect 62 -103 63 -102
rect 67 -103 68 -102
rect 68 -103 69 -102
rect 69 -103 70 -102
rect 70 -103 71 -102
rect 71 -103 72 -102
rect 72 -103 73 -102
rect 73 -103 74 -102
rect 74 -103 75 -102
rect 75 -103 76 -102
rect 76 -103 77 -102
rect 77 -103 78 -102
rect 78 -103 79 -102
rect 79 -103 80 -102
rect 80 -103 81 -102
rect 81 -103 82 -102
rect 82 -103 83 -102
rect 83 -103 84 -102
rect 84 -103 85 -102
rect 85 -103 86 -102
rect 86 -103 87 -102
rect 87 -103 88 -102
rect 88 -103 89 -102
rect 89 -103 90 -102
rect 90 -103 91 -102
rect 91 -103 92 -102
rect 92 -103 93 -102
rect 93 -103 94 -102
rect 94 -103 95 -102
rect 99 -103 100 -102
rect 100 -103 101 -102
rect 101 -103 102 -102
rect 102 -103 103 -102
rect 103 -103 104 -102
rect 104 -103 105 -102
rect 105 -103 106 -102
rect 106 -103 107 -102
rect 107 -103 108 -102
rect 108 -103 109 -102
rect 109 -103 110 -102
rect 110 -103 111 -102
rect 111 -103 112 -102
rect 112 -103 113 -102
rect 113 -103 114 -102
rect 114 -103 115 -102
rect 115 -103 116 -102
rect 116 -103 117 -102
rect 117 -103 118 -102
rect 118 -103 119 -102
rect 119 -103 120 -102
rect 120 -103 121 -102
rect 121 -103 122 -102
rect 122 -103 123 -102
rect 123 -103 124 -102
rect 124 -103 125 -102
rect 125 -103 126 -102
rect 126 -103 127 -102
rect 131 -103 132 -102
rect 132 -103 133 -102
rect 133 -103 134 -102
rect 134 -103 135 -102
rect 135 -103 136 -102
rect 136 -103 137 -102
rect 137 -103 138 -102
rect 138 -103 139 -102
rect 139 -103 140 -102
rect 140 -103 141 -102
rect 141 -103 142 -102
rect 142 -103 143 -102
rect 143 -103 144 -102
rect 144 -103 145 -102
rect 145 -103 146 -102
rect 146 -103 147 -102
rect 147 -103 148 -102
rect 148 -103 149 -102
rect 149 -103 150 -102
rect 150 -103 151 -102
rect 151 -103 152 -102
rect 152 -103 153 -102
rect 153 -103 154 -102
rect 154 -103 155 -102
rect 155 -103 156 -102
rect 156 -103 157 -102
rect 157 -103 158 -102
rect 158 -103 159 -102
rect 163 -103 164 -102
rect 164 -103 165 -102
rect 165 -103 166 -102
rect 166 -103 167 -102
rect 167 -103 168 -102
rect 168 -103 169 -102
rect 169 -103 170 -102
rect 170 -103 171 -102
rect 171 -103 172 -102
rect 172 -103 173 -102
rect 173 -103 174 -102
rect 174 -103 175 -102
rect 175 -103 176 -102
rect 176 -103 177 -102
rect 177 -103 178 -102
rect 178 -103 179 -102
rect 179 -103 180 -102
rect 180 -103 181 -102
rect 181 -103 182 -102
rect 182 -103 183 -102
rect 183 -103 184 -102
rect 184 -103 185 -102
rect 185 -103 186 -102
rect 186 -103 187 -102
rect 187 -103 188 -102
rect 188 -103 189 -102
rect 189 -103 190 -102
rect 190 -103 191 -102
rect 191 -103 192 -102
rect 2 -104 3 -103
rect 3 -104 4 -103
rect 4 -104 5 -103
rect 5 -104 6 -103
rect 6 -104 7 -103
rect 7 -104 8 -103
rect 8 -104 9 -103
rect 9 -104 10 -103
rect 10 -104 11 -103
rect 11 -104 12 -103
rect 12 -104 13 -103
rect 13 -104 14 -103
rect 14 -104 15 -103
rect 15 -104 16 -103
rect 16 -104 17 -103
rect 17 -104 18 -103
rect 18 -104 19 -103
rect 19 -104 20 -103
rect 20 -104 21 -103
rect 21 -104 22 -103
rect 22 -104 23 -103
rect 23 -104 24 -103
rect 24 -104 25 -103
rect 25 -104 26 -103
rect 26 -104 27 -103
rect 27 -104 28 -103
rect 28 -104 29 -103
rect 29 -104 30 -103
rect 30 -104 31 -103
rect 35 -104 36 -103
rect 36 -104 37 -103
rect 37 -104 38 -103
rect 38 -104 39 -103
rect 39 -104 40 -103
rect 40 -104 41 -103
rect 41 -104 42 -103
rect 42 -104 43 -103
rect 43 -104 44 -103
rect 44 -104 45 -103
rect 45 -104 46 -103
rect 46 -104 47 -103
rect 47 -104 48 -103
rect 48 -104 49 -103
rect 49 -104 50 -103
rect 50 -104 51 -103
rect 51 -104 52 -103
rect 52 -104 53 -103
rect 53 -104 54 -103
rect 54 -104 55 -103
rect 55 -104 56 -103
rect 56 -104 57 -103
rect 57 -104 58 -103
rect 58 -104 59 -103
rect 59 -104 60 -103
rect 60 -104 61 -103
rect 61 -104 62 -103
rect 62 -104 63 -103
rect 67 -104 68 -103
rect 68 -104 69 -103
rect 69 -104 70 -103
rect 70 -104 71 -103
rect 71 -104 72 -103
rect 72 -104 73 -103
rect 73 -104 74 -103
rect 74 -104 75 -103
rect 75 -104 76 -103
rect 76 -104 77 -103
rect 77 -104 78 -103
rect 78 -104 79 -103
rect 79 -104 80 -103
rect 80 -104 81 -103
rect 81 -104 82 -103
rect 82 -104 83 -103
rect 83 -104 84 -103
rect 84 -104 85 -103
rect 85 -104 86 -103
rect 86 -104 87 -103
rect 87 -104 88 -103
rect 88 -104 89 -103
rect 89 -104 90 -103
rect 90 -104 91 -103
rect 91 -104 92 -103
rect 92 -104 93 -103
rect 93 -104 94 -103
rect 94 -104 95 -103
rect 99 -104 100 -103
rect 100 -104 101 -103
rect 101 -104 102 -103
rect 102 -104 103 -103
rect 103 -104 104 -103
rect 104 -104 105 -103
rect 105 -104 106 -103
rect 106 -104 107 -103
rect 107 -104 108 -103
rect 108 -104 109 -103
rect 109 -104 110 -103
rect 110 -104 111 -103
rect 111 -104 112 -103
rect 112 -104 113 -103
rect 113 -104 114 -103
rect 114 -104 115 -103
rect 115 -104 116 -103
rect 116 -104 117 -103
rect 117 -104 118 -103
rect 118 -104 119 -103
rect 119 -104 120 -103
rect 120 -104 121 -103
rect 121 -104 122 -103
rect 122 -104 123 -103
rect 123 -104 124 -103
rect 124 -104 125 -103
rect 125 -104 126 -103
rect 126 -104 127 -103
rect 131 -104 132 -103
rect 132 -104 133 -103
rect 133 -104 134 -103
rect 134 -104 135 -103
rect 135 -104 136 -103
rect 136 -104 137 -103
rect 137 -104 138 -103
rect 138 -104 139 -103
rect 139 -104 140 -103
rect 140 -104 141 -103
rect 141 -104 142 -103
rect 142 -104 143 -103
rect 143 -104 144 -103
rect 144 -104 145 -103
rect 145 -104 146 -103
rect 146 -104 147 -103
rect 147 -104 148 -103
rect 148 -104 149 -103
rect 149 -104 150 -103
rect 150 -104 151 -103
rect 151 -104 152 -103
rect 152 -104 153 -103
rect 153 -104 154 -103
rect 154 -104 155 -103
rect 155 -104 156 -103
rect 156 -104 157 -103
rect 157 -104 158 -103
rect 158 -104 159 -103
rect 163 -104 164 -103
rect 164 -104 165 -103
rect 165 -104 166 -103
rect 166 -104 167 -103
rect 167 -104 168 -103
rect 168 -104 169 -103
rect 169 -104 170 -103
rect 170 -104 171 -103
rect 171 -104 172 -103
rect 172 -104 173 -103
rect 173 -104 174 -103
rect 174 -104 175 -103
rect 175 -104 176 -103
rect 176 -104 177 -103
rect 177 -104 178 -103
rect 178 -104 179 -103
rect 179 -104 180 -103
rect 180 -104 181 -103
rect 181 -104 182 -103
rect 182 -104 183 -103
rect 183 -104 184 -103
rect 184 -104 185 -103
rect 185 -104 186 -103
rect 186 -104 187 -103
rect 187 -104 188 -103
rect 188 -104 189 -103
rect 189 -104 190 -103
rect 190 -104 191 -103
rect 191 -104 192 -103
rect 2 -105 3 -104
rect 3 -105 4 -104
rect 4 -105 5 -104
rect 5 -105 6 -104
rect 6 -105 7 -104
rect 7 -105 8 -104
rect 8 -105 9 -104
rect 9 -105 10 -104
rect 10 -105 11 -104
rect 11 -105 12 -104
rect 12 -105 13 -104
rect 13 -105 14 -104
rect 14 -105 15 -104
rect 15 -105 16 -104
rect 16 -105 17 -104
rect 17 -105 18 -104
rect 18 -105 19 -104
rect 19 -105 20 -104
rect 20 -105 21 -104
rect 21 -105 22 -104
rect 22 -105 23 -104
rect 23 -105 24 -104
rect 24 -105 25 -104
rect 25 -105 26 -104
rect 26 -105 27 -104
rect 27 -105 28 -104
rect 28 -105 29 -104
rect 29 -105 30 -104
rect 35 -105 36 -104
rect 36 -105 37 -104
rect 37 -105 38 -104
rect 38 -105 39 -104
rect 39 -105 40 -104
rect 40 -105 41 -104
rect 41 -105 42 -104
rect 42 -105 43 -104
rect 43 -105 44 -104
rect 44 -105 45 -104
rect 45 -105 46 -104
rect 46 -105 47 -104
rect 47 -105 48 -104
rect 48 -105 49 -104
rect 49 -105 50 -104
rect 50 -105 51 -104
rect 51 -105 52 -104
rect 52 -105 53 -104
rect 53 -105 54 -104
rect 54 -105 55 -104
rect 55 -105 56 -104
rect 56 -105 57 -104
rect 57 -105 58 -104
rect 58 -105 59 -104
rect 59 -105 60 -104
rect 60 -105 61 -104
rect 61 -105 62 -104
rect 67 -105 68 -104
rect 68 -105 69 -104
rect 69 -105 70 -104
rect 70 -105 71 -104
rect 71 -105 72 -104
rect 72 -105 73 -104
rect 73 -105 74 -104
rect 74 -105 75 -104
rect 75 -105 76 -104
rect 76 -105 77 -104
rect 77 -105 78 -104
rect 78 -105 79 -104
rect 79 -105 80 -104
rect 80 -105 81 -104
rect 81 -105 82 -104
rect 82 -105 83 -104
rect 83 -105 84 -104
rect 84 -105 85 -104
rect 85 -105 86 -104
rect 86 -105 87 -104
rect 87 -105 88 -104
rect 88 -105 89 -104
rect 89 -105 90 -104
rect 90 -105 91 -104
rect 91 -105 92 -104
rect 92 -105 93 -104
rect 93 -105 94 -104
rect 99 -105 100 -104
rect 100 -105 101 -104
rect 101 -105 102 -104
rect 102 -105 103 -104
rect 103 -105 104 -104
rect 104 -105 105 -104
rect 105 -105 106 -104
rect 106 -105 107 -104
rect 107 -105 108 -104
rect 108 -105 109 -104
rect 109 -105 110 -104
rect 110 -105 111 -104
rect 111 -105 112 -104
rect 112 -105 113 -104
rect 113 -105 114 -104
rect 114 -105 115 -104
rect 115 -105 116 -104
rect 116 -105 117 -104
rect 117 -105 118 -104
rect 118 -105 119 -104
rect 119 -105 120 -104
rect 120 -105 121 -104
rect 121 -105 122 -104
rect 122 -105 123 -104
rect 123 -105 124 -104
rect 124 -105 125 -104
rect 125 -105 126 -104
rect 131 -105 132 -104
rect 132 -105 133 -104
rect 133 -105 134 -104
rect 134 -105 135 -104
rect 135 -105 136 -104
rect 136 -105 137 -104
rect 137 -105 138 -104
rect 138 -105 139 -104
rect 139 -105 140 -104
rect 140 -105 141 -104
rect 141 -105 142 -104
rect 142 -105 143 -104
rect 143 -105 144 -104
rect 144 -105 145 -104
rect 145 -105 146 -104
rect 146 -105 147 -104
rect 147 -105 148 -104
rect 148 -105 149 -104
rect 149 -105 150 -104
rect 150 -105 151 -104
rect 151 -105 152 -104
rect 152 -105 153 -104
rect 153 -105 154 -104
rect 154 -105 155 -104
rect 155 -105 156 -104
rect 156 -105 157 -104
rect 157 -105 158 -104
rect 163 -105 164 -104
rect 164 -105 165 -104
rect 165 -105 166 -104
rect 166 -105 167 -104
rect 167 -105 168 -104
rect 168 -105 169 -104
rect 169 -105 170 -104
rect 170 -105 171 -104
rect 171 -105 172 -104
rect 172 -105 173 -104
rect 173 -105 174 -104
rect 174 -105 175 -104
rect 175 -105 176 -104
rect 176 -105 177 -104
rect 177 -105 178 -104
rect 178 -105 179 -104
rect 179 -105 180 -104
rect 180 -105 181 -104
rect 181 -105 182 -104
rect 182 -105 183 -104
rect 183 -105 184 -104
rect 184 -105 185 -104
rect 185 -105 186 -104
rect 186 -105 187 -104
rect 187 -105 188 -104
rect 188 -105 189 -104
rect 189 -105 190 -104
rect 190 -105 191 -104
rect 191 -105 192 -104
rect 2 -106 3 -105
rect 3 -106 4 -105
rect 4 -106 5 -105
rect 5 -106 6 -105
rect 6 -106 7 -105
rect 7 -106 8 -105
rect 8 -106 9 -105
rect 9 -106 10 -105
rect 10 -106 11 -105
rect 11 -106 12 -105
rect 12 -106 13 -105
rect 13 -106 14 -105
rect 14 -106 15 -105
rect 15 -106 16 -105
rect 16 -106 17 -105
rect 17 -106 18 -105
rect 18 -106 19 -105
rect 19 -106 20 -105
rect 20 -106 21 -105
rect 21 -106 22 -105
rect 22 -106 23 -105
rect 23 -106 24 -105
rect 24 -106 25 -105
rect 41 -106 42 -105
rect 42 -106 43 -105
rect 43 -106 44 -105
rect 44 -106 45 -105
rect 45 -106 46 -105
rect 46 -106 47 -105
rect 47 -106 48 -105
rect 48 -106 49 -105
rect 49 -106 50 -105
rect 50 -106 51 -105
rect 51 -106 52 -105
rect 52 -106 53 -105
rect 53 -106 54 -105
rect 54 -106 55 -105
rect 55 -106 56 -105
rect 56 -106 57 -105
rect 73 -106 74 -105
rect 74 -106 75 -105
rect 75 -106 76 -105
rect 76 -106 77 -105
rect 77 -106 78 -105
rect 78 -106 79 -105
rect 79 -106 80 -105
rect 80 -106 81 -105
rect 81 -106 82 -105
rect 82 -106 83 -105
rect 83 -106 84 -105
rect 84 -106 85 -105
rect 85 -106 86 -105
rect 86 -106 87 -105
rect 87 -106 88 -105
rect 88 -106 89 -105
rect 105 -106 106 -105
rect 106 -106 107 -105
rect 107 -106 108 -105
rect 108 -106 109 -105
rect 109 -106 110 -105
rect 110 -106 111 -105
rect 111 -106 112 -105
rect 112 -106 113 -105
rect 113 -106 114 -105
rect 114 -106 115 -105
rect 115 -106 116 -105
rect 116 -106 117 -105
rect 117 -106 118 -105
rect 118 -106 119 -105
rect 119 -106 120 -105
rect 120 -106 121 -105
rect 137 -106 138 -105
rect 138 -106 139 -105
rect 139 -106 140 -105
rect 140 -106 141 -105
rect 141 -106 142 -105
rect 142 -106 143 -105
rect 143 -106 144 -105
rect 144 -106 145 -105
rect 145 -106 146 -105
rect 146 -106 147 -105
rect 147 -106 148 -105
rect 148 -106 149 -105
rect 149 -106 150 -105
rect 150 -106 151 -105
rect 151 -106 152 -105
rect 152 -106 153 -105
rect 169 -106 170 -105
rect 170 -106 171 -105
rect 171 -106 172 -105
rect 172 -106 173 -105
rect 173 -106 174 -105
rect 174 -106 175 -105
rect 175 -106 176 -105
rect 176 -106 177 -105
rect 177 -106 178 -105
rect 178 -106 179 -105
rect 179 -106 180 -105
rect 180 -106 181 -105
rect 181 -106 182 -105
rect 182 -106 183 -105
rect 183 -106 184 -105
rect 184 -106 185 -105
rect 185 -106 186 -105
rect 186 -106 187 -105
rect 187 -106 188 -105
rect 188 -106 189 -105
rect 189 -106 190 -105
rect 190 -106 191 -105
rect 191 -106 192 -105
rect 2 -107 3 -106
rect 3 -107 4 -106
rect 4 -107 5 -106
rect 5 -107 6 -106
rect 6 -107 7 -106
rect 7 -107 8 -106
rect 8 -107 9 -106
rect 9 -107 10 -106
rect 10 -107 11 -106
rect 11 -107 12 -106
rect 12 -107 13 -106
rect 13 -107 14 -106
rect 14 -107 15 -106
rect 15 -107 16 -106
rect 16 -107 17 -106
rect 17 -107 18 -106
rect 18 -107 19 -106
rect 19 -107 20 -106
rect 20 -107 21 -106
rect 21 -107 22 -106
rect 22 -107 23 -106
rect 23 -107 24 -106
rect 24 -107 25 -106
rect 41 -107 42 -106
rect 42 -107 43 -106
rect 43 -107 44 -106
rect 44 -107 45 -106
rect 45 -107 46 -106
rect 46 -107 47 -106
rect 47 -107 48 -106
rect 48 -107 49 -106
rect 49 -107 50 -106
rect 50 -107 51 -106
rect 51 -107 52 -106
rect 52 -107 53 -106
rect 53 -107 54 -106
rect 54 -107 55 -106
rect 55 -107 56 -106
rect 56 -107 57 -106
rect 73 -107 74 -106
rect 74 -107 75 -106
rect 75 -107 76 -106
rect 76 -107 77 -106
rect 77 -107 78 -106
rect 78 -107 79 -106
rect 79 -107 80 -106
rect 80 -107 81 -106
rect 81 -107 82 -106
rect 82 -107 83 -106
rect 83 -107 84 -106
rect 84 -107 85 -106
rect 85 -107 86 -106
rect 86 -107 87 -106
rect 87 -107 88 -106
rect 88 -107 89 -106
rect 105 -107 106 -106
rect 106 -107 107 -106
rect 107 -107 108 -106
rect 108 -107 109 -106
rect 109 -107 110 -106
rect 110 -107 111 -106
rect 111 -107 112 -106
rect 112 -107 113 -106
rect 113 -107 114 -106
rect 114 -107 115 -106
rect 115 -107 116 -106
rect 116 -107 117 -106
rect 117 -107 118 -106
rect 118 -107 119 -106
rect 119 -107 120 -106
rect 120 -107 121 -106
rect 137 -107 138 -106
rect 138 -107 139 -106
rect 139 -107 140 -106
rect 140 -107 141 -106
rect 141 -107 142 -106
rect 142 -107 143 -106
rect 143 -107 144 -106
rect 144 -107 145 -106
rect 145 -107 146 -106
rect 146 -107 147 -106
rect 147 -107 148 -106
rect 148 -107 149 -106
rect 149 -107 150 -106
rect 150 -107 151 -106
rect 151 -107 152 -106
rect 152 -107 153 -106
rect 169 -107 170 -106
rect 170 -107 171 -106
rect 171 -107 172 -106
rect 172 -107 173 -106
rect 173 -107 174 -106
rect 174 -107 175 -106
rect 175 -107 176 -106
rect 176 -107 177 -106
rect 177 -107 178 -106
rect 178 -107 179 -106
rect 179 -107 180 -106
rect 180 -107 181 -106
rect 181 -107 182 -106
rect 182 -107 183 -106
rect 183 -107 184 -106
rect 184 -107 185 -106
rect 185 -107 186 -106
rect 186 -107 187 -106
rect 187 -107 188 -106
rect 188 -107 189 -106
rect 189 -107 190 -106
rect 190 -107 191 -106
rect 191 -107 192 -106
rect 2 -108 3 -107
rect 3 -108 4 -107
rect 4 -108 5 -107
rect 5 -108 6 -107
rect 6 -108 7 -107
rect 7 -108 8 -107
rect 8 -108 9 -107
rect 9 -108 10 -107
rect 10 -108 11 -107
rect 11 -108 12 -107
rect 12 -108 13 -107
rect 13 -108 14 -107
rect 14 -108 15 -107
rect 15 -108 16 -107
rect 16 -108 17 -107
rect 17 -108 18 -107
rect 18 -108 19 -107
rect 19 -108 20 -107
rect 20 -108 21 -107
rect 21 -108 22 -107
rect 22 -108 23 -107
rect 23 -108 24 -107
rect 24 -108 25 -107
rect 25 -108 26 -107
rect 39 -108 40 -107
rect 40 -108 41 -107
rect 41 -108 42 -107
rect 42 -108 43 -107
rect 43 -108 44 -107
rect 44 -108 45 -107
rect 45 -108 46 -107
rect 46 -108 47 -107
rect 47 -108 48 -107
rect 48 -108 49 -107
rect 49 -108 50 -107
rect 50 -108 51 -107
rect 51 -108 52 -107
rect 52 -108 53 -107
rect 53 -108 54 -107
rect 54 -108 55 -107
rect 55 -108 56 -107
rect 56 -108 57 -107
rect 57 -108 58 -107
rect 71 -108 72 -107
rect 72 -108 73 -107
rect 73 -108 74 -107
rect 74 -108 75 -107
rect 75 -108 76 -107
rect 76 -108 77 -107
rect 77 -108 78 -107
rect 78 -108 79 -107
rect 79 -108 80 -107
rect 80 -108 81 -107
rect 81 -108 82 -107
rect 82 -108 83 -107
rect 83 -108 84 -107
rect 84 -108 85 -107
rect 85 -108 86 -107
rect 86 -108 87 -107
rect 87 -108 88 -107
rect 88 -108 89 -107
rect 89 -108 90 -107
rect 103 -108 104 -107
rect 104 -108 105 -107
rect 105 -108 106 -107
rect 106 -108 107 -107
rect 107 -108 108 -107
rect 108 -108 109 -107
rect 109 -108 110 -107
rect 110 -108 111 -107
rect 111 -108 112 -107
rect 112 -108 113 -107
rect 113 -108 114 -107
rect 114 -108 115 -107
rect 115 -108 116 -107
rect 116 -108 117 -107
rect 117 -108 118 -107
rect 118 -108 119 -107
rect 119 -108 120 -107
rect 120 -108 121 -107
rect 121 -108 122 -107
rect 135 -108 136 -107
rect 136 -108 137 -107
rect 137 -108 138 -107
rect 138 -108 139 -107
rect 139 -108 140 -107
rect 140 -108 141 -107
rect 141 -108 142 -107
rect 142 -108 143 -107
rect 143 -108 144 -107
rect 144 -108 145 -107
rect 145 -108 146 -107
rect 146 -108 147 -107
rect 147 -108 148 -107
rect 148 -108 149 -107
rect 149 -108 150 -107
rect 150 -108 151 -107
rect 151 -108 152 -107
rect 152 -108 153 -107
rect 153 -108 154 -107
rect 167 -108 168 -107
rect 168 -108 169 -107
rect 169 -108 170 -107
rect 170 -108 171 -107
rect 171 -108 172 -107
rect 172 -108 173 -107
rect 173 -108 174 -107
rect 174 -108 175 -107
rect 175 -108 176 -107
rect 176 -108 177 -107
rect 177 -108 178 -107
rect 178 -108 179 -107
rect 179 -108 180 -107
rect 180 -108 181 -107
rect 181 -108 182 -107
rect 182 -108 183 -107
rect 183 -108 184 -107
rect 184 -108 185 -107
rect 185 -108 186 -107
rect 186 -108 187 -107
rect 187 -108 188 -107
rect 188 -108 189 -107
rect 189 -108 190 -107
rect 190 -108 191 -107
rect 191 -108 192 -107
rect 2 -109 3 -108
rect 3 -109 4 -108
rect 4 -109 5 -108
rect 5 -109 6 -108
rect 6 -109 7 -108
rect 7 -109 8 -108
rect 8 -109 9 -108
rect 9 -109 10 -108
rect 10 -109 11 -108
rect 11 -109 12 -108
rect 12 -109 13 -108
rect 13 -109 14 -108
rect 14 -109 15 -108
rect 15 -109 16 -108
rect 16 -109 17 -108
rect 17 -109 18 -108
rect 18 -109 19 -108
rect 19 -109 20 -108
rect 20 -109 21 -108
rect 21 -109 22 -108
rect 22 -109 23 -108
rect 23 -109 24 -108
rect 24 -109 25 -108
rect 25 -109 26 -108
rect 26 -109 27 -108
rect 38 -109 39 -108
rect 39 -109 40 -108
rect 40 -109 41 -108
rect 41 -109 42 -108
rect 42 -109 43 -108
rect 43 -109 44 -108
rect 44 -109 45 -108
rect 45 -109 46 -108
rect 46 -109 47 -108
rect 47 -109 48 -108
rect 48 -109 49 -108
rect 49 -109 50 -108
rect 50 -109 51 -108
rect 51 -109 52 -108
rect 52 -109 53 -108
rect 53 -109 54 -108
rect 54 -109 55 -108
rect 55 -109 56 -108
rect 56 -109 57 -108
rect 57 -109 58 -108
rect 58 -109 59 -108
rect 70 -109 71 -108
rect 71 -109 72 -108
rect 72 -109 73 -108
rect 73 -109 74 -108
rect 74 -109 75 -108
rect 75 -109 76 -108
rect 76 -109 77 -108
rect 77 -109 78 -108
rect 78 -109 79 -108
rect 79 -109 80 -108
rect 80 -109 81 -108
rect 81 -109 82 -108
rect 82 -109 83 -108
rect 83 -109 84 -108
rect 84 -109 85 -108
rect 85 -109 86 -108
rect 86 -109 87 -108
rect 87 -109 88 -108
rect 88 -109 89 -108
rect 89 -109 90 -108
rect 90 -109 91 -108
rect 102 -109 103 -108
rect 103 -109 104 -108
rect 104 -109 105 -108
rect 105 -109 106 -108
rect 106 -109 107 -108
rect 107 -109 108 -108
rect 108 -109 109 -108
rect 109 -109 110 -108
rect 110 -109 111 -108
rect 111 -109 112 -108
rect 112 -109 113 -108
rect 113 -109 114 -108
rect 114 -109 115 -108
rect 115 -109 116 -108
rect 116 -109 117 -108
rect 117 -109 118 -108
rect 118 -109 119 -108
rect 119 -109 120 -108
rect 120 -109 121 -108
rect 121 -109 122 -108
rect 122 -109 123 -108
rect 134 -109 135 -108
rect 135 -109 136 -108
rect 136 -109 137 -108
rect 137 -109 138 -108
rect 138 -109 139 -108
rect 139 -109 140 -108
rect 140 -109 141 -108
rect 141 -109 142 -108
rect 142 -109 143 -108
rect 143 -109 144 -108
rect 144 -109 145 -108
rect 145 -109 146 -108
rect 146 -109 147 -108
rect 147 -109 148 -108
rect 148 -109 149 -108
rect 149 -109 150 -108
rect 150 -109 151 -108
rect 151 -109 152 -108
rect 152 -109 153 -108
rect 153 -109 154 -108
rect 154 -109 155 -108
rect 166 -109 167 -108
rect 167 -109 168 -108
rect 168 -109 169 -108
rect 169 -109 170 -108
rect 170 -109 171 -108
rect 171 -109 172 -108
rect 172 -109 173 -108
rect 173 -109 174 -108
rect 174 -109 175 -108
rect 175 -109 176 -108
rect 176 -109 177 -108
rect 177 -109 178 -108
rect 178 -109 179 -108
rect 179 -109 180 -108
rect 180 -109 181 -108
rect 181 -109 182 -108
rect 182 -109 183 -108
rect 183 -109 184 -108
rect 184 -109 185 -108
rect 185 -109 186 -108
rect 186 -109 187 -108
rect 187 -109 188 -108
rect 188 -109 189 -108
rect 189 -109 190 -108
rect 190 -109 191 -108
rect 191 -109 192 -108
rect 2 -110 3 -109
rect 3 -110 4 -109
rect 4 -110 5 -109
rect 5 -110 6 -109
rect 6 -110 7 -109
rect 7 -110 8 -109
rect 8 -110 9 -109
rect 9 -110 10 -109
rect 10 -110 11 -109
rect 11 -110 12 -109
rect 12 -110 13 -109
rect 13 -110 14 -109
rect 14 -110 15 -109
rect 15 -110 16 -109
rect 16 -110 17 -109
rect 17 -110 18 -109
rect 18 -110 19 -109
rect 19 -110 20 -109
rect 20 -110 21 -109
rect 21 -110 22 -109
rect 22 -110 23 -109
rect 23 -110 24 -109
rect 24 -110 25 -109
rect 25 -110 26 -109
rect 26 -110 27 -109
rect 27 -110 28 -109
rect 37 -110 38 -109
rect 38 -110 39 -109
rect 39 -110 40 -109
rect 40 -110 41 -109
rect 41 -110 42 -109
rect 42 -110 43 -109
rect 43 -110 44 -109
rect 44 -110 45 -109
rect 45 -110 46 -109
rect 46 -110 47 -109
rect 47 -110 48 -109
rect 48 -110 49 -109
rect 49 -110 50 -109
rect 50 -110 51 -109
rect 51 -110 52 -109
rect 52 -110 53 -109
rect 53 -110 54 -109
rect 54 -110 55 -109
rect 55 -110 56 -109
rect 56 -110 57 -109
rect 57 -110 58 -109
rect 58 -110 59 -109
rect 59 -110 60 -109
rect 69 -110 70 -109
rect 70 -110 71 -109
rect 71 -110 72 -109
rect 72 -110 73 -109
rect 73 -110 74 -109
rect 74 -110 75 -109
rect 75 -110 76 -109
rect 76 -110 77 -109
rect 77 -110 78 -109
rect 78 -110 79 -109
rect 79 -110 80 -109
rect 80 -110 81 -109
rect 81 -110 82 -109
rect 82 -110 83 -109
rect 83 -110 84 -109
rect 84 -110 85 -109
rect 85 -110 86 -109
rect 86 -110 87 -109
rect 87 -110 88 -109
rect 88 -110 89 -109
rect 89 -110 90 -109
rect 90 -110 91 -109
rect 91 -110 92 -109
rect 101 -110 102 -109
rect 102 -110 103 -109
rect 103 -110 104 -109
rect 104 -110 105 -109
rect 105 -110 106 -109
rect 106 -110 107 -109
rect 107 -110 108 -109
rect 108 -110 109 -109
rect 109 -110 110 -109
rect 110 -110 111 -109
rect 111 -110 112 -109
rect 112 -110 113 -109
rect 113 -110 114 -109
rect 114 -110 115 -109
rect 115 -110 116 -109
rect 116 -110 117 -109
rect 117 -110 118 -109
rect 118 -110 119 -109
rect 119 -110 120 -109
rect 120 -110 121 -109
rect 121 -110 122 -109
rect 122 -110 123 -109
rect 123 -110 124 -109
rect 133 -110 134 -109
rect 134 -110 135 -109
rect 135 -110 136 -109
rect 136 -110 137 -109
rect 137 -110 138 -109
rect 138 -110 139 -109
rect 139 -110 140 -109
rect 140 -110 141 -109
rect 141 -110 142 -109
rect 142 -110 143 -109
rect 143 -110 144 -109
rect 144 -110 145 -109
rect 145 -110 146 -109
rect 146 -110 147 -109
rect 147 -110 148 -109
rect 148 -110 149 -109
rect 149 -110 150 -109
rect 150 -110 151 -109
rect 151 -110 152 -109
rect 152 -110 153 -109
rect 153 -110 154 -109
rect 154 -110 155 -109
rect 155 -110 156 -109
rect 165 -110 166 -109
rect 166 -110 167 -109
rect 167 -110 168 -109
rect 168 -110 169 -109
rect 169 -110 170 -109
rect 170 -110 171 -109
rect 171 -110 172 -109
rect 172 -110 173 -109
rect 173 -110 174 -109
rect 174 -110 175 -109
rect 175 -110 176 -109
rect 176 -110 177 -109
rect 177 -110 178 -109
rect 178 -110 179 -109
rect 179 -110 180 -109
rect 180 -110 181 -109
rect 181 -110 182 -109
rect 182 -110 183 -109
rect 183 -110 184 -109
rect 184 -110 185 -109
rect 185 -110 186 -109
rect 186 -110 187 -109
rect 187 -110 188 -109
rect 188 -110 189 -109
rect 189 -110 190 -109
rect 190 -110 191 -109
rect 191 -110 192 -109
rect 2 -111 3 -110
rect 3 -111 4 -110
rect 4 -111 5 -110
rect 5 -111 6 -110
rect 6 -111 7 -110
rect 7 -111 8 -110
rect 8 -111 9 -110
rect 9 -111 10 -110
rect 10 -111 11 -110
rect 11 -111 12 -110
rect 12 -111 13 -110
rect 13 -111 14 -110
rect 14 -111 15 -110
rect 15 -111 16 -110
rect 16 -111 17 -110
rect 17 -111 18 -110
rect 18 -111 19 -110
rect 19 -111 20 -110
rect 20 -111 21 -110
rect 21 -111 22 -110
rect 22 -111 23 -110
rect 23 -111 24 -110
rect 24 -111 25 -110
rect 25 -111 26 -110
rect 26 -111 27 -110
rect 27 -111 28 -110
rect 37 -111 38 -110
rect 38 -111 39 -110
rect 39 -111 40 -110
rect 40 -111 41 -110
rect 41 -111 42 -110
rect 42 -111 43 -110
rect 43 -111 44 -110
rect 44 -111 45 -110
rect 45 -111 46 -110
rect 46 -111 47 -110
rect 47 -111 48 -110
rect 48 -111 49 -110
rect 49 -111 50 -110
rect 50 -111 51 -110
rect 51 -111 52 -110
rect 52 -111 53 -110
rect 53 -111 54 -110
rect 54 -111 55 -110
rect 55 -111 56 -110
rect 56 -111 57 -110
rect 57 -111 58 -110
rect 58 -111 59 -110
rect 59 -111 60 -110
rect 69 -111 70 -110
rect 70 -111 71 -110
rect 71 -111 72 -110
rect 72 -111 73 -110
rect 73 -111 74 -110
rect 74 -111 75 -110
rect 75 -111 76 -110
rect 76 -111 77 -110
rect 77 -111 78 -110
rect 78 -111 79 -110
rect 79 -111 80 -110
rect 80 -111 81 -110
rect 81 -111 82 -110
rect 82 -111 83 -110
rect 83 -111 84 -110
rect 84 -111 85 -110
rect 85 -111 86 -110
rect 86 -111 87 -110
rect 87 -111 88 -110
rect 88 -111 89 -110
rect 89 -111 90 -110
rect 90 -111 91 -110
rect 91 -111 92 -110
rect 101 -111 102 -110
rect 102 -111 103 -110
rect 103 -111 104 -110
rect 104 -111 105 -110
rect 105 -111 106 -110
rect 106 -111 107 -110
rect 107 -111 108 -110
rect 108 -111 109 -110
rect 109 -111 110 -110
rect 110 -111 111 -110
rect 111 -111 112 -110
rect 112 -111 113 -110
rect 113 -111 114 -110
rect 114 -111 115 -110
rect 115 -111 116 -110
rect 116 -111 117 -110
rect 117 -111 118 -110
rect 118 -111 119 -110
rect 119 -111 120 -110
rect 120 -111 121 -110
rect 121 -111 122 -110
rect 122 -111 123 -110
rect 123 -111 124 -110
rect 133 -111 134 -110
rect 134 -111 135 -110
rect 135 -111 136 -110
rect 136 -111 137 -110
rect 137 -111 138 -110
rect 138 -111 139 -110
rect 139 -111 140 -110
rect 140 -111 141 -110
rect 141 -111 142 -110
rect 142 -111 143 -110
rect 143 -111 144 -110
rect 144 -111 145 -110
rect 145 -111 146 -110
rect 146 -111 147 -110
rect 147 -111 148 -110
rect 148 -111 149 -110
rect 149 -111 150 -110
rect 150 -111 151 -110
rect 151 -111 152 -110
rect 152 -111 153 -110
rect 153 -111 154 -110
rect 154 -111 155 -110
rect 155 -111 156 -110
rect 165 -111 166 -110
rect 166 -111 167 -110
rect 167 -111 168 -110
rect 168 -111 169 -110
rect 169 -111 170 -110
rect 170 -111 171 -110
rect 171 -111 172 -110
rect 172 -111 173 -110
rect 173 -111 174 -110
rect 174 -111 175 -110
rect 175 -111 176 -110
rect 176 -111 177 -110
rect 177 -111 178 -110
rect 178 -111 179 -110
rect 179 -111 180 -110
rect 180 -111 181 -110
rect 181 -111 182 -110
rect 182 -111 183 -110
rect 183 -111 184 -110
rect 184 -111 185 -110
rect 185 -111 186 -110
rect 186 -111 187 -110
rect 187 -111 188 -110
rect 188 -111 189 -110
rect 189 -111 190 -110
rect 190 -111 191 -110
rect 191 -111 192 -110
rect 2 -112 3 -111
rect 3 -112 4 -111
rect 4 -112 5 -111
rect 5 -112 6 -111
rect 6 -112 7 -111
rect 7 -112 8 -111
rect 8 -112 9 -111
rect 9 -112 10 -111
rect 10 -112 11 -111
rect 11 -112 12 -111
rect 12 -112 13 -111
rect 13 -112 14 -111
rect 14 -112 15 -111
rect 15 -112 16 -111
rect 16 -112 17 -111
rect 17 -112 18 -111
rect 18 -112 19 -111
rect 19 -112 20 -111
rect 20 -112 21 -111
rect 21 -112 22 -111
rect 22 -112 23 -111
rect 23 -112 24 -111
rect 24 -112 25 -111
rect 25 -112 26 -111
rect 26 -112 27 -111
rect 27 -112 28 -111
rect 37 -112 38 -111
rect 38 -112 39 -111
rect 39 -112 40 -111
rect 40 -112 41 -111
rect 41 -112 42 -111
rect 42 -112 43 -111
rect 43 -112 44 -111
rect 44 -112 45 -111
rect 45 -112 46 -111
rect 46 -112 47 -111
rect 47 -112 48 -111
rect 48 -112 49 -111
rect 49 -112 50 -111
rect 50 -112 51 -111
rect 51 -112 52 -111
rect 52 -112 53 -111
rect 53 -112 54 -111
rect 54 -112 55 -111
rect 55 -112 56 -111
rect 56 -112 57 -111
rect 57 -112 58 -111
rect 58 -112 59 -111
rect 59 -112 60 -111
rect 69 -112 70 -111
rect 70 -112 71 -111
rect 71 -112 72 -111
rect 72 -112 73 -111
rect 73 -112 74 -111
rect 74 -112 75 -111
rect 75 -112 76 -111
rect 76 -112 77 -111
rect 77 -112 78 -111
rect 78 -112 79 -111
rect 79 -112 80 -111
rect 80 -112 81 -111
rect 81 -112 82 -111
rect 82 -112 83 -111
rect 83 -112 84 -111
rect 84 -112 85 -111
rect 85 -112 86 -111
rect 86 -112 87 -111
rect 87 -112 88 -111
rect 88 -112 89 -111
rect 89 -112 90 -111
rect 90 -112 91 -111
rect 91 -112 92 -111
rect 101 -112 102 -111
rect 102 -112 103 -111
rect 103 -112 104 -111
rect 104 -112 105 -111
rect 105 -112 106 -111
rect 106 -112 107 -111
rect 107 -112 108 -111
rect 108 -112 109 -111
rect 109 -112 110 -111
rect 110 -112 111 -111
rect 111 -112 112 -111
rect 112 -112 113 -111
rect 113 -112 114 -111
rect 114 -112 115 -111
rect 115 -112 116 -111
rect 116 -112 117 -111
rect 117 -112 118 -111
rect 118 -112 119 -111
rect 119 -112 120 -111
rect 120 -112 121 -111
rect 121 -112 122 -111
rect 122 -112 123 -111
rect 123 -112 124 -111
rect 133 -112 134 -111
rect 134 -112 135 -111
rect 135 -112 136 -111
rect 136 -112 137 -111
rect 137 -112 138 -111
rect 138 -112 139 -111
rect 139 -112 140 -111
rect 140 -112 141 -111
rect 141 -112 142 -111
rect 142 -112 143 -111
rect 143 -112 144 -111
rect 144 -112 145 -111
rect 145 -112 146 -111
rect 146 -112 147 -111
rect 147 -112 148 -111
rect 148 -112 149 -111
rect 149 -112 150 -111
rect 150 -112 151 -111
rect 151 -112 152 -111
rect 152 -112 153 -111
rect 153 -112 154 -111
rect 154 -112 155 -111
rect 155 -112 156 -111
rect 165 -112 166 -111
rect 166 -112 167 -111
rect 167 -112 168 -111
rect 168 -112 169 -111
rect 169 -112 170 -111
rect 170 -112 171 -111
rect 171 -112 172 -111
rect 172 -112 173 -111
rect 173 -112 174 -111
rect 174 -112 175 -111
rect 175 -112 176 -111
rect 176 -112 177 -111
rect 177 -112 178 -111
rect 178 -112 179 -111
rect 179 -112 180 -111
rect 180 -112 181 -111
rect 181 -112 182 -111
rect 182 -112 183 -111
rect 183 -112 184 -111
rect 184 -112 185 -111
rect 185 -112 186 -111
rect 186 -112 187 -111
rect 187 -112 188 -111
rect 188 -112 189 -111
rect 189 -112 190 -111
rect 190 -112 191 -111
rect 191 -112 192 -111
rect 2 -113 3 -112
rect 3 -113 4 -112
rect 4 -113 5 -112
rect 5 -113 6 -112
rect 6 -113 7 -112
rect 7 -113 8 -112
rect 8 -113 9 -112
rect 9 -113 10 -112
rect 10 -113 11 -112
rect 11 -113 12 -112
rect 12 -113 13 -112
rect 13 -113 14 -112
rect 14 -113 15 -112
rect 15 -113 16 -112
rect 16 -113 17 -112
rect 17 -113 18 -112
rect 18 -113 19 -112
rect 19 -113 20 -112
rect 20 -113 21 -112
rect 21 -113 22 -112
rect 22 -113 23 -112
rect 23 -113 24 -112
rect 24 -113 25 -112
rect 25 -113 26 -112
rect 26 -113 27 -112
rect 27 -113 28 -112
rect 32 -113 33 -112
rect 38 -113 39 -112
rect 39 -113 40 -112
rect 40 -113 41 -112
rect 41 -113 42 -112
rect 42 -113 43 -112
rect 43 -113 44 -112
rect 44 -113 45 -112
rect 45 -113 46 -112
rect 46 -113 47 -112
rect 47 -113 48 -112
rect 48 -113 49 -112
rect 49 -113 50 -112
rect 50 -113 51 -112
rect 51 -113 52 -112
rect 52 -113 53 -112
rect 53 -113 54 -112
rect 54 -113 55 -112
rect 55 -113 56 -112
rect 56 -113 57 -112
rect 57 -113 58 -112
rect 58 -113 59 -112
rect 59 -113 60 -112
rect 64 -113 65 -112
rect 70 -113 71 -112
rect 71 -113 72 -112
rect 72 -113 73 -112
rect 73 -113 74 -112
rect 74 -113 75 -112
rect 75 -113 76 -112
rect 76 -113 77 -112
rect 77 -113 78 -112
rect 78 -113 79 -112
rect 79 -113 80 -112
rect 80 -113 81 -112
rect 81 -113 82 -112
rect 82 -113 83 -112
rect 83 -113 84 -112
rect 84 -113 85 -112
rect 85 -113 86 -112
rect 86 -113 87 -112
rect 87 -113 88 -112
rect 88 -113 89 -112
rect 89 -113 90 -112
rect 90 -113 91 -112
rect 91 -113 92 -112
rect 96 -113 97 -112
rect 102 -113 103 -112
rect 103 -113 104 -112
rect 104 -113 105 -112
rect 105 -113 106 -112
rect 106 -113 107 -112
rect 107 -113 108 -112
rect 108 -113 109 -112
rect 109 -113 110 -112
rect 110 -113 111 -112
rect 111 -113 112 -112
rect 112 -113 113 -112
rect 113 -113 114 -112
rect 114 -113 115 -112
rect 115 -113 116 -112
rect 116 -113 117 -112
rect 117 -113 118 -112
rect 118 -113 119 -112
rect 119 -113 120 -112
rect 120 -113 121 -112
rect 121 -113 122 -112
rect 122 -113 123 -112
rect 123 -113 124 -112
rect 128 -113 129 -112
rect 134 -113 135 -112
rect 135 -113 136 -112
rect 136 -113 137 -112
rect 137 -113 138 -112
rect 138 -113 139 -112
rect 139 -113 140 -112
rect 140 -113 141 -112
rect 141 -113 142 -112
rect 142 -113 143 -112
rect 143 -113 144 -112
rect 144 -113 145 -112
rect 145 -113 146 -112
rect 146 -113 147 -112
rect 147 -113 148 -112
rect 148 -113 149 -112
rect 149 -113 150 -112
rect 150 -113 151 -112
rect 151 -113 152 -112
rect 152 -113 153 -112
rect 153 -113 154 -112
rect 154 -113 155 -112
rect 155 -113 156 -112
rect 160 -113 161 -112
rect 166 -113 167 -112
rect 167 -113 168 -112
rect 168 -113 169 -112
rect 169 -113 170 -112
rect 170 -113 171 -112
rect 171 -113 172 -112
rect 172 -113 173 -112
rect 173 -113 174 -112
rect 174 -113 175 -112
rect 175 -113 176 -112
rect 176 -113 177 -112
rect 177 -113 178 -112
rect 178 -113 179 -112
rect 179 -113 180 -112
rect 180 -113 181 -112
rect 181 -113 182 -112
rect 182 -113 183 -112
rect 183 -113 184 -112
rect 184 -113 185 -112
rect 185 -113 186 -112
rect 186 -113 187 -112
rect 187 -113 188 -112
rect 188 -113 189 -112
rect 189 -113 190 -112
rect 190 -113 191 -112
rect 191 -113 192 -112
rect 2 -114 3 -113
rect 3 -114 4 -113
rect 4 -114 5 -113
rect 5 -114 6 -113
rect 6 -114 7 -113
rect 7 -114 8 -113
rect 8 -114 9 -113
rect 9 -114 10 -113
rect 10 -114 11 -113
rect 11 -114 12 -113
rect 12 -114 13 -113
rect 13 -114 14 -113
rect 14 -114 15 -113
rect 15 -114 16 -113
rect 16 -114 17 -113
rect 17 -114 18 -113
rect 18 -114 19 -113
rect 19 -114 20 -113
rect 20 -114 21 -113
rect 21 -114 22 -113
rect 22 -114 23 -113
rect 23 -114 24 -113
rect 24 -114 25 -113
rect 25 -114 26 -113
rect 26 -114 27 -113
rect 27 -114 28 -113
rect 31 -114 32 -113
rect 32 -114 33 -113
rect 33 -114 34 -113
rect 38 -114 39 -113
rect 39 -114 40 -113
rect 40 -114 41 -113
rect 41 -114 42 -113
rect 42 -114 43 -113
rect 43 -114 44 -113
rect 44 -114 45 -113
rect 45 -114 46 -113
rect 46 -114 47 -113
rect 47 -114 48 -113
rect 48 -114 49 -113
rect 49 -114 50 -113
rect 50 -114 51 -113
rect 51 -114 52 -113
rect 52 -114 53 -113
rect 53 -114 54 -113
rect 54 -114 55 -113
rect 55 -114 56 -113
rect 56 -114 57 -113
rect 57 -114 58 -113
rect 58 -114 59 -113
rect 59 -114 60 -113
rect 63 -114 64 -113
rect 64 -114 65 -113
rect 65 -114 66 -113
rect 70 -114 71 -113
rect 71 -114 72 -113
rect 72 -114 73 -113
rect 73 -114 74 -113
rect 74 -114 75 -113
rect 75 -114 76 -113
rect 76 -114 77 -113
rect 77 -114 78 -113
rect 78 -114 79 -113
rect 79 -114 80 -113
rect 80 -114 81 -113
rect 81 -114 82 -113
rect 82 -114 83 -113
rect 83 -114 84 -113
rect 84 -114 85 -113
rect 85 -114 86 -113
rect 86 -114 87 -113
rect 87 -114 88 -113
rect 88 -114 89 -113
rect 89 -114 90 -113
rect 90 -114 91 -113
rect 91 -114 92 -113
rect 95 -114 96 -113
rect 96 -114 97 -113
rect 97 -114 98 -113
rect 102 -114 103 -113
rect 103 -114 104 -113
rect 104 -114 105 -113
rect 105 -114 106 -113
rect 106 -114 107 -113
rect 107 -114 108 -113
rect 108 -114 109 -113
rect 109 -114 110 -113
rect 110 -114 111 -113
rect 111 -114 112 -113
rect 112 -114 113 -113
rect 113 -114 114 -113
rect 114 -114 115 -113
rect 115 -114 116 -113
rect 116 -114 117 -113
rect 117 -114 118 -113
rect 118 -114 119 -113
rect 119 -114 120 -113
rect 120 -114 121 -113
rect 121 -114 122 -113
rect 122 -114 123 -113
rect 123 -114 124 -113
rect 127 -114 128 -113
rect 128 -114 129 -113
rect 129 -114 130 -113
rect 134 -114 135 -113
rect 135 -114 136 -113
rect 136 -114 137 -113
rect 137 -114 138 -113
rect 138 -114 139 -113
rect 139 -114 140 -113
rect 140 -114 141 -113
rect 141 -114 142 -113
rect 142 -114 143 -113
rect 143 -114 144 -113
rect 144 -114 145 -113
rect 145 -114 146 -113
rect 146 -114 147 -113
rect 147 -114 148 -113
rect 148 -114 149 -113
rect 149 -114 150 -113
rect 150 -114 151 -113
rect 151 -114 152 -113
rect 152 -114 153 -113
rect 153 -114 154 -113
rect 154 -114 155 -113
rect 155 -114 156 -113
rect 159 -114 160 -113
rect 160 -114 161 -113
rect 161 -114 162 -113
rect 166 -114 167 -113
rect 167 -114 168 -113
rect 168 -114 169 -113
rect 169 -114 170 -113
rect 170 -114 171 -113
rect 171 -114 172 -113
rect 172 -114 173 -113
rect 173 -114 174 -113
rect 174 -114 175 -113
rect 175 -114 176 -113
rect 176 -114 177 -113
rect 177 -114 178 -113
rect 178 -114 179 -113
rect 179 -114 180 -113
rect 180 -114 181 -113
rect 181 -114 182 -113
rect 182 -114 183 -113
rect 183 -114 184 -113
rect 184 -114 185 -113
rect 185 -114 186 -113
rect 186 -114 187 -113
rect 187 -114 188 -113
rect 188 -114 189 -113
rect 189 -114 190 -113
rect 190 -114 191 -113
rect 191 -114 192 -113
rect 2 -115 3 -114
rect 3 -115 4 -114
rect 4 -115 5 -114
rect 5 -115 6 -114
rect 6 -115 7 -114
rect 7 -115 8 -114
rect 8 -115 9 -114
rect 9 -115 10 -114
rect 10 -115 11 -114
rect 11 -115 12 -114
rect 12 -115 13 -114
rect 13 -115 14 -114
rect 14 -115 15 -114
rect 18 -115 19 -114
rect 19 -115 20 -114
rect 20 -115 21 -114
rect 21 -115 22 -114
rect 22 -115 23 -114
rect 23 -115 24 -114
rect 24 -115 25 -114
rect 25 -115 26 -114
rect 26 -115 27 -114
rect 27 -115 28 -114
rect 30 -115 31 -114
rect 31 -115 32 -114
rect 32 -115 33 -114
rect 33 -115 34 -114
rect 34 -115 35 -114
rect 38 -115 39 -114
rect 39 -115 40 -114
rect 40 -115 41 -114
rect 41 -115 42 -114
rect 42 -115 43 -114
rect 43 -115 44 -114
rect 44 -115 45 -114
rect 45 -115 46 -114
rect 46 -115 47 -114
rect 50 -115 51 -114
rect 51 -115 52 -114
rect 52 -115 53 -114
rect 53 -115 54 -114
rect 54 -115 55 -114
rect 55 -115 56 -114
rect 56 -115 57 -114
rect 57 -115 58 -114
rect 58 -115 59 -114
rect 59 -115 60 -114
rect 62 -115 63 -114
rect 63 -115 64 -114
rect 64 -115 65 -114
rect 65 -115 66 -114
rect 66 -115 67 -114
rect 70 -115 71 -114
rect 71 -115 72 -114
rect 72 -115 73 -114
rect 73 -115 74 -114
rect 74 -115 75 -114
rect 75 -115 76 -114
rect 76 -115 77 -114
rect 77 -115 78 -114
rect 78 -115 79 -114
rect 82 -115 83 -114
rect 83 -115 84 -114
rect 84 -115 85 -114
rect 85 -115 86 -114
rect 86 -115 87 -114
rect 87 -115 88 -114
rect 88 -115 89 -114
rect 89 -115 90 -114
rect 90 -115 91 -114
rect 91 -115 92 -114
rect 94 -115 95 -114
rect 95 -115 96 -114
rect 96 -115 97 -114
rect 97 -115 98 -114
rect 98 -115 99 -114
rect 102 -115 103 -114
rect 103 -115 104 -114
rect 104 -115 105 -114
rect 105 -115 106 -114
rect 106 -115 107 -114
rect 107 -115 108 -114
rect 108 -115 109 -114
rect 109 -115 110 -114
rect 110 -115 111 -114
rect 114 -115 115 -114
rect 115 -115 116 -114
rect 116 -115 117 -114
rect 117 -115 118 -114
rect 118 -115 119 -114
rect 119 -115 120 -114
rect 120 -115 121 -114
rect 121 -115 122 -114
rect 122 -115 123 -114
rect 123 -115 124 -114
rect 126 -115 127 -114
rect 127 -115 128 -114
rect 128 -115 129 -114
rect 129 -115 130 -114
rect 130 -115 131 -114
rect 134 -115 135 -114
rect 135 -115 136 -114
rect 136 -115 137 -114
rect 137 -115 138 -114
rect 138 -115 139 -114
rect 139 -115 140 -114
rect 140 -115 141 -114
rect 141 -115 142 -114
rect 142 -115 143 -114
rect 146 -115 147 -114
rect 147 -115 148 -114
rect 148 -115 149 -114
rect 149 -115 150 -114
rect 150 -115 151 -114
rect 151 -115 152 -114
rect 152 -115 153 -114
rect 153 -115 154 -114
rect 154 -115 155 -114
rect 155 -115 156 -114
rect 158 -115 159 -114
rect 159 -115 160 -114
rect 160 -115 161 -114
rect 161 -115 162 -114
rect 162 -115 163 -114
rect 166 -115 167 -114
rect 167 -115 168 -114
rect 168 -115 169 -114
rect 169 -115 170 -114
rect 170 -115 171 -114
rect 171 -115 172 -114
rect 172 -115 173 -114
rect 173 -115 174 -114
rect 174 -115 175 -114
rect 178 -115 179 -114
rect 179 -115 180 -114
rect 180 -115 181 -114
rect 181 -115 182 -114
rect 182 -115 183 -114
rect 183 -115 184 -114
rect 184 -115 185 -114
rect 185 -115 186 -114
rect 186 -115 187 -114
rect 187 -115 188 -114
rect 188 -115 189 -114
rect 189 -115 190 -114
rect 190 -115 191 -114
rect 191 -115 192 -114
rect 2 -116 3 -115
rect 3 -116 4 -115
rect 4 -116 5 -115
rect 5 -116 6 -115
rect 6 -116 7 -115
rect 7 -116 8 -115
rect 8 -116 9 -115
rect 9 -116 10 -115
rect 10 -116 11 -115
rect 11 -116 12 -115
rect 12 -116 13 -115
rect 13 -116 14 -115
rect 14 -116 15 -115
rect 18 -116 19 -115
rect 19 -116 20 -115
rect 20 -116 21 -115
rect 21 -116 22 -115
rect 22 -116 23 -115
rect 23 -116 24 -115
rect 24 -116 25 -115
rect 25 -116 26 -115
rect 26 -116 27 -115
rect 27 -116 28 -115
rect 28 -116 29 -115
rect 29 -116 30 -115
rect 30 -116 31 -115
rect 31 -116 32 -115
rect 32 -116 33 -115
rect 33 -116 34 -115
rect 34 -116 35 -115
rect 35 -116 36 -115
rect 36 -116 37 -115
rect 37 -116 38 -115
rect 38 -116 39 -115
rect 39 -116 40 -115
rect 40 -116 41 -115
rect 41 -116 42 -115
rect 42 -116 43 -115
rect 43 -116 44 -115
rect 44 -116 45 -115
rect 45 -116 46 -115
rect 46 -116 47 -115
rect 50 -116 51 -115
rect 51 -116 52 -115
rect 52 -116 53 -115
rect 53 -116 54 -115
rect 54 -116 55 -115
rect 55 -116 56 -115
rect 56 -116 57 -115
rect 57 -116 58 -115
rect 58 -116 59 -115
rect 59 -116 60 -115
rect 60 -116 61 -115
rect 61 -116 62 -115
rect 62 -116 63 -115
rect 63 -116 64 -115
rect 64 -116 65 -115
rect 65 -116 66 -115
rect 66 -116 67 -115
rect 67 -116 68 -115
rect 68 -116 69 -115
rect 69 -116 70 -115
rect 70 -116 71 -115
rect 71 -116 72 -115
rect 72 -116 73 -115
rect 73 -116 74 -115
rect 74 -116 75 -115
rect 75 -116 76 -115
rect 76 -116 77 -115
rect 77 -116 78 -115
rect 78 -116 79 -115
rect 82 -116 83 -115
rect 83 -116 84 -115
rect 84 -116 85 -115
rect 85 -116 86 -115
rect 86 -116 87 -115
rect 87 -116 88 -115
rect 88 -116 89 -115
rect 89 -116 90 -115
rect 90 -116 91 -115
rect 91 -116 92 -115
rect 92 -116 93 -115
rect 93 -116 94 -115
rect 94 -116 95 -115
rect 95 -116 96 -115
rect 96 -116 97 -115
rect 97 -116 98 -115
rect 98 -116 99 -115
rect 99 -116 100 -115
rect 100 -116 101 -115
rect 101 -116 102 -115
rect 102 -116 103 -115
rect 103 -116 104 -115
rect 104 -116 105 -115
rect 105 -116 106 -115
rect 106 -116 107 -115
rect 107 -116 108 -115
rect 108 -116 109 -115
rect 109 -116 110 -115
rect 110 -116 111 -115
rect 114 -116 115 -115
rect 115 -116 116 -115
rect 116 -116 117 -115
rect 117 -116 118 -115
rect 118 -116 119 -115
rect 119 -116 120 -115
rect 120 -116 121 -115
rect 121 -116 122 -115
rect 122 -116 123 -115
rect 123 -116 124 -115
rect 124 -116 125 -115
rect 125 -116 126 -115
rect 126 -116 127 -115
rect 127 -116 128 -115
rect 128 -116 129 -115
rect 129 -116 130 -115
rect 130 -116 131 -115
rect 131 -116 132 -115
rect 132 -116 133 -115
rect 133 -116 134 -115
rect 134 -116 135 -115
rect 135 -116 136 -115
rect 136 -116 137 -115
rect 137 -116 138 -115
rect 138 -116 139 -115
rect 139 -116 140 -115
rect 140 -116 141 -115
rect 141 -116 142 -115
rect 142 -116 143 -115
rect 146 -116 147 -115
rect 147 -116 148 -115
rect 148 -116 149 -115
rect 149 -116 150 -115
rect 150 -116 151 -115
rect 151 -116 152 -115
rect 152 -116 153 -115
rect 153 -116 154 -115
rect 154 -116 155 -115
rect 155 -116 156 -115
rect 156 -116 157 -115
rect 157 -116 158 -115
rect 158 -116 159 -115
rect 159 -116 160 -115
rect 160 -116 161 -115
rect 161 -116 162 -115
rect 162 -116 163 -115
rect 163 -116 164 -115
rect 164 -116 165 -115
rect 165 -116 166 -115
rect 166 -116 167 -115
rect 167 -116 168 -115
rect 168 -116 169 -115
rect 169 -116 170 -115
rect 170 -116 171 -115
rect 171 -116 172 -115
rect 172 -116 173 -115
rect 173 -116 174 -115
rect 174 -116 175 -115
rect 178 -116 179 -115
rect 179 -116 180 -115
rect 180 -116 181 -115
rect 181 -116 182 -115
rect 182 -116 183 -115
rect 183 -116 184 -115
rect 184 -116 185 -115
rect 185 -116 186 -115
rect 186 -116 187 -115
rect 187 -116 188 -115
rect 188 -116 189 -115
rect 189 -116 190 -115
rect 190 -116 191 -115
rect 191 -116 192 -115
rect 2 -117 3 -116
rect 3 -117 4 -116
rect 4 -117 5 -116
rect 5 -117 6 -116
rect 6 -117 7 -116
rect 7 -117 8 -116
rect 8 -117 9 -116
rect 9 -117 10 -116
rect 10 -117 11 -116
rect 11 -117 12 -116
rect 12 -117 13 -116
rect 13 -117 14 -116
rect 14 -117 15 -116
rect 19 -117 20 -116
rect 20 -117 21 -116
rect 21 -117 22 -116
rect 22 -117 23 -116
rect 23 -117 24 -116
rect 24 -117 25 -116
rect 25 -117 26 -116
rect 26 -117 27 -116
rect 27 -117 28 -116
rect 28 -117 29 -116
rect 29 -117 30 -116
rect 30 -117 31 -116
rect 31 -117 32 -116
rect 32 -117 33 -116
rect 33 -117 34 -116
rect 34 -117 35 -116
rect 35 -117 36 -116
rect 36 -117 37 -116
rect 37 -117 38 -116
rect 38 -117 39 -116
rect 39 -117 40 -116
rect 40 -117 41 -116
rect 41 -117 42 -116
rect 42 -117 43 -116
rect 43 -117 44 -116
rect 44 -117 45 -116
rect 45 -117 46 -116
rect 46 -117 47 -116
rect 51 -117 52 -116
rect 52 -117 53 -116
rect 53 -117 54 -116
rect 54 -117 55 -116
rect 55 -117 56 -116
rect 56 -117 57 -116
rect 57 -117 58 -116
rect 58 -117 59 -116
rect 59 -117 60 -116
rect 60 -117 61 -116
rect 61 -117 62 -116
rect 62 -117 63 -116
rect 63 -117 64 -116
rect 64 -117 65 -116
rect 65 -117 66 -116
rect 66 -117 67 -116
rect 67 -117 68 -116
rect 68 -117 69 -116
rect 69 -117 70 -116
rect 70 -117 71 -116
rect 71 -117 72 -116
rect 72 -117 73 -116
rect 73 -117 74 -116
rect 74 -117 75 -116
rect 75 -117 76 -116
rect 76 -117 77 -116
rect 77 -117 78 -116
rect 78 -117 79 -116
rect 83 -117 84 -116
rect 84 -117 85 -116
rect 85 -117 86 -116
rect 86 -117 87 -116
rect 87 -117 88 -116
rect 88 -117 89 -116
rect 89 -117 90 -116
rect 90 -117 91 -116
rect 91 -117 92 -116
rect 92 -117 93 -116
rect 93 -117 94 -116
rect 94 -117 95 -116
rect 95 -117 96 -116
rect 96 -117 97 -116
rect 97 -117 98 -116
rect 98 -117 99 -116
rect 99 -117 100 -116
rect 100 -117 101 -116
rect 101 -117 102 -116
rect 102 -117 103 -116
rect 103 -117 104 -116
rect 104 -117 105 -116
rect 105 -117 106 -116
rect 106 -117 107 -116
rect 107 -117 108 -116
rect 108 -117 109 -116
rect 109 -117 110 -116
rect 110 -117 111 -116
rect 115 -117 116 -116
rect 116 -117 117 -116
rect 117 -117 118 -116
rect 118 -117 119 -116
rect 119 -117 120 -116
rect 120 -117 121 -116
rect 121 -117 122 -116
rect 122 -117 123 -116
rect 123 -117 124 -116
rect 124 -117 125 -116
rect 125 -117 126 -116
rect 126 -117 127 -116
rect 127 -117 128 -116
rect 128 -117 129 -116
rect 129 -117 130 -116
rect 130 -117 131 -116
rect 131 -117 132 -116
rect 132 -117 133 -116
rect 133 -117 134 -116
rect 134 -117 135 -116
rect 135 -117 136 -116
rect 136 -117 137 -116
rect 137 -117 138 -116
rect 138 -117 139 -116
rect 139 -117 140 -116
rect 140 -117 141 -116
rect 141 -117 142 -116
rect 142 -117 143 -116
rect 147 -117 148 -116
rect 148 -117 149 -116
rect 149 -117 150 -116
rect 150 -117 151 -116
rect 151 -117 152 -116
rect 152 -117 153 -116
rect 153 -117 154 -116
rect 154 -117 155 -116
rect 155 -117 156 -116
rect 156 -117 157 -116
rect 157 -117 158 -116
rect 158 -117 159 -116
rect 159 -117 160 -116
rect 160 -117 161 -116
rect 161 -117 162 -116
rect 162 -117 163 -116
rect 163 -117 164 -116
rect 164 -117 165 -116
rect 165 -117 166 -116
rect 166 -117 167 -116
rect 167 -117 168 -116
rect 168 -117 169 -116
rect 169 -117 170 -116
rect 170 -117 171 -116
rect 171 -117 172 -116
rect 172 -117 173 -116
rect 173 -117 174 -116
rect 174 -117 175 -116
rect 179 -117 180 -116
rect 180 -117 181 -116
rect 181 -117 182 -116
rect 182 -117 183 -116
rect 183 -117 184 -116
rect 184 -117 185 -116
rect 185 -117 186 -116
rect 186 -117 187 -116
rect 187 -117 188 -116
rect 188 -117 189 -116
rect 189 -117 190 -116
rect 190 -117 191 -116
rect 191 -117 192 -116
rect 2 -118 3 -117
rect 3 -118 4 -117
rect 4 -118 5 -117
rect 5 -118 6 -117
rect 6 -118 7 -117
rect 7 -118 8 -117
rect 8 -118 9 -117
rect 9 -118 10 -117
rect 10 -118 11 -117
rect 11 -118 12 -117
rect 12 -118 13 -117
rect 13 -118 14 -117
rect 14 -118 15 -117
rect 19 -118 20 -117
rect 20 -118 21 -117
rect 21 -118 22 -117
rect 22 -118 23 -117
rect 23 -118 24 -117
rect 24 -118 25 -117
rect 25 -118 26 -117
rect 26 -118 27 -117
rect 27 -118 28 -117
rect 28 -118 29 -117
rect 29 -118 30 -117
rect 30 -118 31 -117
rect 31 -118 32 -117
rect 32 -118 33 -117
rect 33 -118 34 -117
rect 34 -118 35 -117
rect 35 -118 36 -117
rect 36 -118 37 -117
rect 37 -118 38 -117
rect 38 -118 39 -117
rect 39 -118 40 -117
rect 40 -118 41 -117
rect 41 -118 42 -117
rect 42 -118 43 -117
rect 43 -118 44 -117
rect 44 -118 45 -117
rect 45 -118 46 -117
rect 46 -118 47 -117
rect 51 -118 52 -117
rect 52 -118 53 -117
rect 53 -118 54 -117
rect 54 -118 55 -117
rect 55 -118 56 -117
rect 56 -118 57 -117
rect 57 -118 58 -117
rect 58 -118 59 -117
rect 59 -118 60 -117
rect 60 -118 61 -117
rect 61 -118 62 -117
rect 62 -118 63 -117
rect 63 -118 64 -117
rect 64 -118 65 -117
rect 65 -118 66 -117
rect 66 -118 67 -117
rect 67 -118 68 -117
rect 68 -118 69 -117
rect 69 -118 70 -117
rect 70 -118 71 -117
rect 71 -118 72 -117
rect 72 -118 73 -117
rect 73 -118 74 -117
rect 74 -118 75 -117
rect 75 -118 76 -117
rect 76 -118 77 -117
rect 77 -118 78 -117
rect 78 -118 79 -117
rect 83 -118 84 -117
rect 84 -118 85 -117
rect 85 -118 86 -117
rect 86 -118 87 -117
rect 87 -118 88 -117
rect 88 -118 89 -117
rect 89 -118 90 -117
rect 90 -118 91 -117
rect 91 -118 92 -117
rect 92 -118 93 -117
rect 93 -118 94 -117
rect 94 -118 95 -117
rect 95 -118 96 -117
rect 96 -118 97 -117
rect 97 -118 98 -117
rect 98 -118 99 -117
rect 99 -118 100 -117
rect 100 -118 101 -117
rect 101 -118 102 -117
rect 102 -118 103 -117
rect 103 -118 104 -117
rect 104 -118 105 -117
rect 105 -118 106 -117
rect 106 -118 107 -117
rect 107 -118 108 -117
rect 108 -118 109 -117
rect 109 -118 110 -117
rect 110 -118 111 -117
rect 115 -118 116 -117
rect 116 -118 117 -117
rect 117 -118 118 -117
rect 118 -118 119 -117
rect 119 -118 120 -117
rect 120 -118 121 -117
rect 121 -118 122 -117
rect 122 -118 123 -117
rect 123 -118 124 -117
rect 124 -118 125 -117
rect 125 -118 126 -117
rect 126 -118 127 -117
rect 127 -118 128 -117
rect 128 -118 129 -117
rect 129 -118 130 -117
rect 130 -118 131 -117
rect 131 -118 132 -117
rect 132 -118 133 -117
rect 133 -118 134 -117
rect 134 -118 135 -117
rect 135 -118 136 -117
rect 136 -118 137 -117
rect 137 -118 138 -117
rect 138 -118 139 -117
rect 139 -118 140 -117
rect 140 -118 141 -117
rect 141 -118 142 -117
rect 142 -118 143 -117
rect 147 -118 148 -117
rect 148 -118 149 -117
rect 149 -118 150 -117
rect 150 -118 151 -117
rect 151 -118 152 -117
rect 152 -118 153 -117
rect 153 -118 154 -117
rect 154 -118 155 -117
rect 155 -118 156 -117
rect 156 -118 157 -117
rect 157 -118 158 -117
rect 158 -118 159 -117
rect 159 -118 160 -117
rect 160 -118 161 -117
rect 161 -118 162 -117
rect 162 -118 163 -117
rect 163 -118 164 -117
rect 164 -118 165 -117
rect 165 -118 166 -117
rect 166 -118 167 -117
rect 167 -118 168 -117
rect 168 -118 169 -117
rect 169 -118 170 -117
rect 170 -118 171 -117
rect 171 -118 172 -117
rect 172 -118 173 -117
rect 173 -118 174 -117
rect 174 -118 175 -117
rect 179 -118 180 -117
rect 180 -118 181 -117
rect 181 -118 182 -117
rect 182 -118 183 -117
rect 183 -118 184 -117
rect 184 -118 185 -117
rect 185 -118 186 -117
rect 186 -118 187 -117
rect 187 -118 188 -117
rect 188 -118 189 -117
rect 189 -118 190 -117
rect 190 -118 191 -117
rect 191 -118 192 -117
rect 192 -118 193 -117
rect 193 -118 194 -117
rect 194 -118 195 -117
rect 195 -118 196 -117
rect 196 -118 197 -117
rect 197 -118 198 -117
rect 198 -118 199 -117
rect 199 -118 200 -117
rect 200 -118 201 -117
rect 201 -118 202 -117
rect 202 -118 203 -117
rect 203 -118 204 -117
rect 204 -118 205 -117
rect 205 -118 206 -117
rect 206 -118 207 -117
rect 207 -118 208 -117
rect 208 -118 209 -117
rect 209 -118 210 -117
rect 210 -118 211 -117
rect 211 -118 212 -117
rect 212 -118 213 -117
rect 213 -118 214 -117
rect 214 -118 215 -117
rect 215 -118 216 -117
rect 216 -118 217 -117
rect 217 -118 218 -117
rect 218 -118 219 -117
rect 219 -118 220 -117
rect 220 -118 221 -117
rect 221 -118 222 -117
rect 222 -118 223 -117
rect 223 -118 224 -117
rect 224 -118 225 -117
rect 225 -118 226 -117
rect 226 -118 227 -117
rect 227 -118 228 -117
rect 228 -118 229 -117
rect 229 -118 230 -117
rect 230 -118 231 -117
rect 231 -118 232 -117
rect 232 -118 233 -117
rect 233 -118 234 -117
rect 234 -118 235 -117
rect 235 -118 236 -117
rect 236 -118 237 -117
rect 237 -118 238 -117
rect 238 -118 239 -117
rect 239 -118 240 -117
rect 240 -118 241 -117
rect 241 -118 242 -117
rect 242 -118 243 -117
rect 243 -118 244 -117
rect 244 -118 245 -117
rect 245 -118 246 -117
rect 246 -118 247 -117
rect 247 -118 248 -117
rect 248 -118 249 -117
rect 249 -118 250 -117
rect 250 -118 251 -117
rect 251 -118 252 -117
rect 252 -118 253 -117
rect 253 -118 254 -117
rect 254 -118 255 -117
rect 255 -118 256 -117
rect 256 -118 257 -117
rect 257 -118 258 -117
rect 258 -118 259 -117
rect 259 -118 260 -117
rect 260 -118 261 -117
rect 261 -118 262 -117
rect 262 -118 263 -117
rect 263 -118 264 -117
rect 264 -118 265 -117
rect 265 -118 266 -117
rect 266 -118 267 -117
rect 267 -118 268 -117
rect 268 -118 269 -117
rect 269 -118 270 -117
rect 270 -118 271 -117
rect 271 -118 272 -117
rect 272 -118 273 -117
rect 273 -118 274 -117
rect 274 -118 275 -117
rect 275 -118 276 -117
rect 276 -118 277 -117
rect 277 -118 278 -117
rect 278 -118 279 -117
rect 279 -118 280 -117
rect 280 -118 281 -117
rect 281 -118 282 -117
rect 282 -118 283 -117
rect 283 -118 284 -117
rect 284 -118 285 -117
rect 285 -118 286 -117
rect 286 -118 287 -117
rect 287 -118 288 -117
rect 288 -118 289 -117
rect 289 -118 290 -117
rect 290 -118 291 -117
rect 291 -118 292 -117
rect 292 -118 293 -117
rect 293 -118 294 -117
rect 294 -118 295 -117
rect 295 -118 296 -117
rect 296 -118 297 -117
rect 297 -118 298 -117
rect 298 -118 299 -117
rect 299 -118 300 -117
rect 300 -118 301 -117
rect 301 -118 302 -117
rect 302 -118 303 -117
rect 303 -118 304 -117
rect 304 -118 305 -117
rect 305 -118 306 -117
rect 306 -118 307 -117
rect 307 -118 308 -117
rect 308 -118 309 -117
rect 309 -118 310 -117
rect 310 -118 311 -117
rect 311 -118 312 -117
rect 312 -118 313 -117
rect 313 -118 314 -117
rect 314 -118 315 -117
rect 315 -118 316 -117
rect 316 -118 317 -117
rect 317 -118 318 -117
rect 318 -118 319 -117
rect 319 -118 320 -117
rect 320 -118 321 -117
rect 321 -118 322 -117
rect 322 -118 323 -117
rect 323 -118 324 -117
rect 324 -118 325 -117
rect 325 -118 326 -117
rect 326 -118 327 -117
rect 327 -118 328 -117
rect 328 -118 329 -117
rect 329 -118 330 -117
rect 330 -118 331 -117
rect 331 -118 332 -117
rect 332 -118 333 -117
rect 333 -118 334 -117
rect 334 -118 335 -117
rect 335 -118 336 -117
rect 336 -118 337 -117
rect 337 -118 338 -117
rect 338 -118 339 -117
rect 339 -118 340 -117
rect 340 -118 341 -117
rect 341 -118 342 -117
rect 342 -118 343 -117
rect 343 -118 344 -117
rect 344 -118 345 -117
rect 345 -118 346 -117
rect 346 -118 347 -117
rect 347 -118 348 -117
rect 348 -118 349 -117
rect 349 -118 350 -117
rect 350 -118 351 -117
rect 351 -118 352 -117
rect 352 -118 353 -117
rect 353 -118 354 -117
rect 354 -118 355 -117
rect 355 -118 356 -117
rect 356 -118 357 -117
rect 357 -118 358 -117
rect 358 -118 359 -117
rect 359 -118 360 -117
rect 360 -118 361 -117
rect 361 -118 362 -117
rect 362 -118 363 -117
rect 363 -118 364 -117
rect 364 -118 365 -117
rect 365 -118 366 -117
rect 366 -118 367 -117
rect 367 -118 368 -117
rect 368 -118 369 -117
rect 369 -118 370 -117
rect 370 -118 371 -117
rect 371 -118 372 -117
rect 372 -118 373 -117
rect 373 -118 374 -117
rect 374 -118 375 -117
rect 375 -118 376 -117
rect 376 -118 377 -117
rect 377 -118 378 -117
rect 378 -118 379 -117
rect 379 -118 380 -117
rect 380 -118 381 -117
rect 381 -118 382 -117
rect 382 -118 383 -117
rect 383 -118 384 -117
rect 384 -118 385 -117
rect 385 -118 386 -117
rect 386 -118 387 -117
rect 387 -118 388 -117
rect 388 -118 389 -117
rect 389 -118 390 -117
rect 390 -118 391 -117
rect 391 -118 392 -117
rect 392 -118 393 -117
rect 393 -118 394 -117
rect 394 -118 395 -117
rect 395 -118 396 -117
rect 396 -118 397 -117
rect 397 -118 398 -117
rect 398 -118 399 -117
rect 399 -118 400 -117
rect 400 -118 401 -117
rect 401 -118 402 -117
rect 402 -118 403 -117
rect 403 -118 404 -117
rect 404 -118 405 -117
rect 405 -118 406 -117
rect 406 -118 407 -117
rect 407 -118 408 -117
rect 408 -118 409 -117
rect 409 -118 410 -117
rect 410 -118 411 -117
rect 411 -118 412 -117
rect 412 -118 413 -117
rect 413 -118 414 -117
rect 414 -118 415 -117
rect 415 -118 416 -117
rect 416 -118 417 -117
rect 417 -118 418 -117
rect 418 -118 419 -117
rect 419 -118 420 -117
rect 420 -118 421 -117
rect 421 -118 422 -117
rect 422 -118 423 -117
rect 423 -118 424 -117
rect 424 -118 425 -117
rect 425 -118 426 -117
rect 426 -118 427 -117
rect 427 -118 428 -117
rect 428 -118 429 -117
rect 429 -118 430 -117
rect 430 -118 431 -117
rect 431 -118 432 -117
rect 432 -118 433 -117
rect 433 -118 434 -117
rect 434 -118 435 -117
rect 435 -118 436 -117
rect 436 -118 437 -117
rect 437 -118 438 -117
rect 438 -118 439 -117
rect 439 -118 440 -117
rect 440 -118 441 -117
rect 441 -118 442 -117
rect 442 -118 443 -117
rect 443 -118 444 -117
rect 444 -118 445 -117
rect 445 -118 446 -117
rect 446 -118 447 -117
rect 447 -118 448 -117
rect 448 -118 449 -117
rect 449 -118 450 -117
rect 450 -118 451 -117
rect 451 -118 452 -117
rect 452 -118 453 -117
rect 453 -118 454 -117
rect 454 -118 455 -117
rect 455 -118 456 -117
rect 456 -118 457 -117
rect 457 -118 458 -117
rect 458 -118 459 -117
rect 459 -118 460 -117
rect 460 -118 461 -117
rect 461 -118 462 -117
rect 462 -118 463 -117
rect 463 -118 464 -117
rect 464 -118 465 -117
rect 465 -118 466 -117
rect 466 -118 467 -117
rect 467 -118 468 -117
rect 468 -118 469 -117
rect 469 -118 470 -117
rect 470 -118 471 -117
rect 471 -118 472 -117
rect 472 -118 473 -117
rect 473 -118 474 -117
rect 474 -118 475 -117
rect 475 -118 476 -117
rect 476 -118 477 -117
rect 477 -118 478 -117
rect 478 -118 479 -117
rect 479 -118 480 -117
rect 2 -119 3 -118
rect 3 -119 4 -118
rect 4 -119 5 -118
rect 5 -119 6 -118
rect 6 -119 7 -118
rect 7 -119 8 -118
rect 8 -119 9 -118
rect 25 -119 26 -118
rect 26 -119 27 -118
rect 27 -119 28 -118
rect 28 -119 29 -118
rect 29 -119 30 -118
rect 30 -119 31 -118
rect 31 -119 32 -118
rect 32 -119 33 -118
rect 33 -119 34 -118
rect 34 -119 35 -118
rect 35 -119 36 -118
rect 36 -119 37 -118
rect 37 -119 38 -118
rect 38 -119 39 -118
rect 39 -119 40 -118
rect 40 -119 41 -118
rect 57 -119 58 -118
rect 58 -119 59 -118
rect 59 -119 60 -118
rect 60 -119 61 -118
rect 61 -119 62 -118
rect 62 -119 63 -118
rect 63 -119 64 -118
rect 64 -119 65 -118
rect 65 -119 66 -118
rect 66 -119 67 -118
rect 67 -119 68 -118
rect 68 -119 69 -118
rect 69 -119 70 -118
rect 70 -119 71 -118
rect 71 -119 72 -118
rect 72 -119 73 -118
rect 89 -119 90 -118
rect 90 -119 91 -118
rect 91 -119 92 -118
rect 92 -119 93 -118
rect 93 -119 94 -118
rect 94 -119 95 -118
rect 95 -119 96 -118
rect 96 -119 97 -118
rect 97 -119 98 -118
rect 98 -119 99 -118
rect 99 -119 100 -118
rect 100 -119 101 -118
rect 101 -119 102 -118
rect 102 -119 103 -118
rect 103 -119 104 -118
rect 104 -119 105 -118
rect 121 -119 122 -118
rect 122 -119 123 -118
rect 123 -119 124 -118
rect 124 -119 125 -118
rect 125 -119 126 -118
rect 126 -119 127 -118
rect 127 -119 128 -118
rect 128 -119 129 -118
rect 129 -119 130 -118
rect 130 -119 131 -118
rect 131 -119 132 -118
rect 132 -119 133 -118
rect 133 -119 134 -118
rect 134 -119 135 -118
rect 135 -119 136 -118
rect 136 -119 137 -118
rect 153 -119 154 -118
rect 154 -119 155 -118
rect 155 -119 156 -118
rect 156 -119 157 -118
rect 157 -119 158 -118
rect 158 -119 159 -118
rect 159 -119 160 -118
rect 160 -119 161 -118
rect 161 -119 162 -118
rect 162 -119 163 -118
rect 163 -119 164 -118
rect 164 -119 165 -118
rect 165 -119 166 -118
rect 166 -119 167 -118
rect 167 -119 168 -118
rect 168 -119 169 -118
rect 185 -119 186 -118
rect 186 -119 187 -118
rect 187 -119 188 -118
rect 188 -119 189 -118
rect 189 -119 190 -118
rect 190 -119 191 -118
rect 191 -119 192 -118
rect 192 -119 193 -118
rect 193 -119 194 -118
rect 194 -119 195 -118
rect 195 -119 196 -118
rect 196 -119 197 -118
rect 197 -119 198 -118
rect 198 -119 199 -118
rect 199 -119 200 -118
rect 200 -119 201 -118
rect 201 -119 202 -118
rect 202 -119 203 -118
rect 203 -119 204 -118
rect 204 -119 205 -118
rect 205 -119 206 -118
rect 206 -119 207 -118
rect 207 -119 208 -118
rect 208 -119 209 -118
rect 209 -119 210 -118
rect 210 -119 211 -118
rect 211 -119 212 -118
rect 212 -119 213 -118
rect 213 -119 214 -118
rect 214 -119 215 -118
rect 215 -119 216 -118
rect 216 -119 217 -118
rect 217 -119 218 -118
rect 218 -119 219 -118
rect 219 -119 220 -118
rect 220 -119 221 -118
rect 221 -119 222 -118
rect 222 -119 223 -118
rect 223 -119 224 -118
rect 224 -119 225 -118
rect 225 -119 226 -118
rect 226 -119 227 -118
rect 227 -119 228 -118
rect 228 -119 229 -118
rect 229 -119 230 -118
rect 230 -119 231 -118
rect 231 -119 232 -118
rect 232 -119 233 -118
rect 233 -119 234 -118
rect 234 -119 235 -118
rect 235 -119 236 -118
rect 236 -119 237 -118
rect 237 -119 238 -118
rect 238 -119 239 -118
rect 239 -119 240 -118
rect 240 -119 241 -118
rect 241 -119 242 -118
rect 242 -119 243 -118
rect 243 -119 244 -118
rect 244 -119 245 -118
rect 245 -119 246 -118
rect 246 -119 247 -118
rect 247 -119 248 -118
rect 248 -119 249 -118
rect 249 -119 250 -118
rect 250 -119 251 -118
rect 251 -119 252 -118
rect 252 -119 253 -118
rect 253 -119 254 -118
rect 254 -119 255 -118
rect 255 -119 256 -118
rect 256 -119 257 -118
rect 257 -119 258 -118
rect 258 -119 259 -118
rect 259 -119 260 -118
rect 260 -119 261 -118
rect 261 -119 262 -118
rect 262 -119 263 -118
rect 263 -119 264 -118
rect 264 -119 265 -118
rect 265 -119 266 -118
rect 266 -119 267 -118
rect 267 -119 268 -118
rect 268 -119 269 -118
rect 269 -119 270 -118
rect 270 -119 271 -118
rect 271 -119 272 -118
rect 272 -119 273 -118
rect 273 -119 274 -118
rect 274 -119 275 -118
rect 275 -119 276 -118
rect 276 -119 277 -118
rect 277 -119 278 -118
rect 278 -119 279 -118
rect 279 -119 280 -118
rect 280 -119 281 -118
rect 281 -119 282 -118
rect 282 -119 283 -118
rect 283 -119 284 -118
rect 284 -119 285 -118
rect 285 -119 286 -118
rect 286 -119 287 -118
rect 287 -119 288 -118
rect 288 -119 289 -118
rect 289 -119 290 -118
rect 290 -119 291 -118
rect 291 -119 292 -118
rect 292 -119 293 -118
rect 293 -119 294 -118
rect 294 -119 295 -118
rect 295 -119 296 -118
rect 296 -119 297 -118
rect 297 -119 298 -118
rect 298 -119 299 -118
rect 299 -119 300 -118
rect 300 -119 301 -118
rect 301 -119 302 -118
rect 302 -119 303 -118
rect 303 -119 304 -118
rect 304 -119 305 -118
rect 305 -119 306 -118
rect 306 -119 307 -118
rect 307 -119 308 -118
rect 308 -119 309 -118
rect 309 -119 310 -118
rect 310 -119 311 -118
rect 311 -119 312 -118
rect 312 -119 313 -118
rect 313 -119 314 -118
rect 314 -119 315 -118
rect 315 -119 316 -118
rect 316 -119 317 -118
rect 317 -119 318 -118
rect 318 -119 319 -118
rect 319 -119 320 -118
rect 320 -119 321 -118
rect 321 -119 322 -118
rect 322 -119 323 -118
rect 323 -119 324 -118
rect 324 -119 325 -118
rect 325 -119 326 -118
rect 326 -119 327 -118
rect 327 -119 328 -118
rect 328 -119 329 -118
rect 329 -119 330 -118
rect 330 -119 331 -118
rect 331 -119 332 -118
rect 332 -119 333 -118
rect 333 -119 334 -118
rect 334 -119 335 -118
rect 335 -119 336 -118
rect 336 -119 337 -118
rect 337 -119 338 -118
rect 338 -119 339 -118
rect 339 -119 340 -118
rect 340 -119 341 -118
rect 341 -119 342 -118
rect 342 -119 343 -118
rect 343 -119 344 -118
rect 344 -119 345 -118
rect 345 -119 346 -118
rect 346 -119 347 -118
rect 347 -119 348 -118
rect 348 -119 349 -118
rect 349 -119 350 -118
rect 350 -119 351 -118
rect 351 -119 352 -118
rect 352 -119 353 -118
rect 353 -119 354 -118
rect 354 -119 355 -118
rect 355 -119 356 -118
rect 356 -119 357 -118
rect 357 -119 358 -118
rect 358 -119 359 -118
rect 359 -119 360 -118
rect 360 -119 361 -118
rect 361 -119 362 -118
rect 362 -119 363 -118
rect 363 -119 364 -118
rect 364 -119 365 -118
rect 365 -119 366 -118
rect 366 -119 367 -118
rect 367 -119 368 -118
rect 368 -119 369 -118
rect 369 -119 370 -118
rect 370 -119 371 -118
rect 371 -119 372 -118
rect 372 -119 373 -118
rect 373 -119 374 -118
rect 374 -119 375 -118
rect 375 -119 376 -118
rect 376 -119 377 -118
rect 377 -119 378 -118
rect 378 -119 379 -118
rect 379 -119 380 -118
rect 380 -119 381 -118
rect 381 -119 382 -118
rect 382 -119 383 -118
rect 383 -119 384 -118
rect 384 -119 385 -118
rect 385 -119 386 -118
rect 386 -119 387 -118
rect 387 -119 388 -118
rect 388 -119 389 -118
rect 389 -119 390 -118
rect 390 -119 391 -118
rect 391 -119 392 -118
rect 392 -119 393 -118
rect 393 -119 394 -118
rect 394 -119 395 -118
rect 395 -119 396 -118
rect 396 -119 397 -118
rect 397 -119 398 -118
rect 398 -119 399 -118
rect 399 -119 400 -118
rect 400 -119 401 -118
rect 401 -119 402 -118
rect 402 -119 403 -118
rect 403 -119 404 -118
rect 404 -119 405 -118
rect 405 -119 406 -118
rect 406 -119 407 -118
rect 407 -119 408 -118
rect 408 -119 409 -118
rect 409 -119 410 -118
rect 410 -119 411 -118
rect 411 -119 412 -118
rect 412 -119 413 -118
rect 413 -119 414 -118
rect 414 -119 415 -118
rect 415 -119 416 -118
rect 416 -119 417 -118
rect 417 -119 418 -118
rect 418 -119 419 -118
rect 419 -119 420 -118
rect 420 -119 421 -118
rect 421 -119 422 -118
rect 422 -119 423 -118
rect 423 -119 424 -118
rect 424 -119 425 -118
rect 425 -119 426 -118
rect 426 -119 427 -118
rect 427 -119 428 -118
rect 428 -119 429 -118
rect 429 -119 430 -118
rect 430 -119 431 -118
rect 431 -119 432 -118
rect 432 -119 433 -118
rect 433 -119 434 -118
rect 434 -119 435 -118
rect 435 -119 436 -118
rect 436 -119 437 -118
rect 437 -119 438 -118
rect 438 -119 439 -118
rect 439 -119 440 -118
rect 440 -119 441 -118
rect 441 -119 442 -118
rect 442 -119 443 -118
rect 443 -119 444 -118
rect 444 -119 445 -118
rect 445 -119 446 -118
rect 446 -119 447 -118
rect 447 -119 448 -118
rect 448 -119 449 -118
rect 449 -119 450 -118
rect 450 -119 451 -118
rect 451 -119 452 -118
rect 452 -119 453 -118
rect 453 -119 454 -118
rect 454 -119 455 -118
rect 455 -119 456 -118
rect 456 -119 457 -118
rect 457 -119 458 -118
rect 458 -119 459 -118
rect 459 -119 460 -118
rect 460 -119 461 -118
rect 461 -119 462 -118
rect 462 -119 463 -118
rect 463 -119 464 -118
rect 464 -119 465 -118
rect 465 -119 466 -118
rect 466 -119 467 -118
rect 467 -119 468 -118
rect 468 -119 469 -118
rect 469 -119 470 -118
rect 470 -119 471 -118
rect 471 -119 472 -118
rect 472 -119 473 -118
rect 473 -119 474 -118
rect 474 -119 475 -118
rect 475 -119 476 -118
rect 476 -119 477 -118
rect 477 -119 478 -118
rect 478 -119 479 -118
rect 479 -119 480 -118
rect 2 -120 3 -119
rect 3 -120 4 -119
rect 4 -120 5 -119
rect 5 -120 6 -119
rect 6 -120 7 -119
rect 7 -120 8 -119
rect 8 -120 9 -119
rect 25 -120 26 -119
rect 26 -120 27 -119
rect 27 -120 28 -119
rect 28 -120 29 -119
rect 29 -120 30 -119
rect 30 -120 31 -119
rect 31 -120 32 -119
rect 32 -120 33 -119
rect 33 -120 34 -119
rect 34 -120 35 -119
rect 35 -120 36 -119
rect 36 -120 37 -119
rect 37 -120 38 -119
rect 38 -120 39 -119
rect 39 -120 40 -119
rect 40 -120 41 -119
rect 57 -120 58 -119
rect 58 -120 59 -119
rect 59 -120 60 -119
rect 60 -120 61 -119
rect 61 -120 62 -119
rect 62 -120 63 -119
rect 63 -120 64 -119
rect 64 -120 65 -119
rect 65 -120 66 -119
rect 66 -120 67 -119
rect 67 -120 68 -119
rect 68 -120 69 -119
rect 69 -120 70 -119
rect 70 -120 71 -119
rect 71 -120 72 -119
rect 72 -120 73 -119
rect 89 -120 90 -119
rect 90 -120 91 -119
rect 91 -120 92 -119
rect 92 -120 93 -119
rect 93 -120 94 -119
rect 94 -120 95 -119
rect 95 -120 96 -119
rect 96 -120 97 -119
rect 97 -120 98 -119
rect 98 -120 99 -119
rect 99 -120 100 -119
rect 100 -120 101 -119
rect 101 -120 102 -119
rect 102 -120 103 -119
rect 103 -120 104 -119
rect 104 -120 105 -119
rect 121 -120 122 -119
rect 122 -120 123 -119
rect 123 -120 124 -119
rect 124 -120 125 -119
rect 125 -120 126 -119
rect 126 -120 127 -119
rect 127 -120 128 -119
rect 128 -120 129 -119
rect 129 -120 130 -119
rect 130 -120 131 -119
rect 131 -120 132 -119
rect 132 -120 133 -119
rect 133 -120 134 -119
rect 134 -120 135 -119
rect 135 -120 136 -119
rect 136 -120 137 -119
rect 153 -120 154 -119
rect 154 -120 155 -119
rect 155 -120 156 -119
rect 156 -120 157 -119
rect 157 -120 158 -119
rect 158 -120 159 -119
rect 159 -120 160 -119
rect 160 -120 161 -119
rect 161 -120 162 -119
rect 162 -120 163 -119
rect 163 -120 164 -119
rect 164 -120 165 -119
rect 165 -120 166 -119
rect 166 -120 167 -119
rect 167 -120 168 -119
rect 168 -120 169 -119
rect 185 -120 186 -119
rect 186 -120 187 -119
rect 187 -120 188 -119
rect 188 -120 189 -119
rect 189 -120 190 -119
rect 190 -120 191 -119
rect 191 -120 192 -119
rect 192 -120 193 -119
rect 193 -120 194 -119
rect 194 -120 195 -119
rect 195 -120 196 -119
rect 196 -120 197 -119
rect 197 -120 198 -119
rect 198 -120 199 -119
rect 199 -120 200 -119
rect 200 -120 201 -119
rect 201 -120 202 -119
rect 202 -120 203 -119
rect 203 -120 204 -119
rect 204 -120 205 -119
rect 205 -120 206 -119
rect 206 -120 207 -119
rect 207 -120 208 -119
rect 208 -120 209 -119
rect 209 -120 210 -119
rect 210 -120 211 -119
rect 211 -120 212 -119
rect 212 -120 213 -119
rect 213 -120 214 -119
rect 214 -120 215 -119
rect 215 -120 216 -119
rect 216 -120 217 -119
rect 217 -120 218 -119
rect 218 -120 219 -119
rect 219 -120 220 -119
rect 220 -120 221 -119
rect 221 -120 222 -119
rect 222 -120 223 -119
rect 223 -120 224 -119
rect 224 -120 225 -119
rect 225 -120 226 -119
rect 226 -120 227 -119
rect 227 -120 228 -119
rect 228 -120 229 -119
rect 229 -120 230 -119
rect 230 -120 231 -119
rect 231 -120 232 -119
rect 232 -120 233 -119
rect 233 -120 234 -119
rect 234 -120 235 -119
rect 235 -120 236 -119
rect 236 -120 237 -119
rect 237 -120 238 -119
rect 238 -120 239 -119
rect 239 -120 240 -119
rect 240 -120 241 -119
rect 241 -120 242 -119
rect 242 -120 243 -119
rect 243 -120 244 -119
rect 244 -120 245 -119
rect 245 -120 246 -119
rect 246 -120 247 -119
rect 247 -120 248 -119
rect 248 -120 249 -119
rect 249 -120 250 -119
rect 250 -120 251 -119
rect 251 -120 252 -119
rect 252 -120 253 -119
rect 253 -120 254 -119
rect 254 -120 255 -119
rect 255 -120 256 -119
rect 256 -120 257 -119
rect 257 -120 258 -119
rect 258 -120 259 -119
rect 259 -120 260 -119
rect 260 -120 261 -119
rect 261 -120 262 -119
rect 262 -120 263 -119
rect 263 -120 264 -119
rect 264 -120 265 -119
rect 265 -120 266 -119
rect 266 -120 267 -119
rect 267 -120 268 -119
rect 268 -120 269 -119
rect 269 -120 270 -119
rect 270 -120 271 -119
rect 271 -120 272 -119
rect 272 -120 273 -119
rect 273 -120 274 -119
rect 274 -120 275 -119
rect 275 -120 276 -119
rect 276 -120 277 -119
rect 277 -120 278 -119
rect 278 -120 279 -119
rect 279 -120 280 -119
rect 280 -120 281 -119
rect 281 -120 282 -119
rect 282 -120 283 -119
rect 283 -120 284 -119
rect 284 -120 285 -119
rect 285 -120 286 -119
rect 286 -120 287 -119
rect 287 -120 288 -119
rect 288 -120 289 -119
rect 289 -120 290 -119
rect 290 -120 291 -119
rect 291 -120 292 -119
rect 292 -120 293 -119
rect 293 -120 294 -119
rect 294 -120 295 -119
rect 295 -120 296 -119
rect 296 -120 297 -119
rect 297 -120 298 -119
rect 298 -120 299 -119
rect 299 -120 300 -119
rect 300 -120 301 -119
rect 301 -120 302 -119
rect 302 -120 303 -119
rect 303 -120 304 -119
rect 304 -120 305 -119
rect 305 -120 306 -119
rect 306 -120 307 -119
rect 307 -120 308 -119
rect 308 -120 309 -119
rect 309 -120 310 -119
rect 310 -120 311 -119
rect 311 -120 312 -119
rect 312 -120 313 -119
rect 313 -120 314 -119
rect 314 -120 315 -119
rect 315 -120 316 -119
rect 316 -120 317 -119
rect 317 -120 318 -119
rect 318 -120 319 -119
rect 319 -120 320 -119
rect 320 -120 321 -119
rect 321 -120 322 -119
rect 322 -120 323 -119
rect 323 -120 324 -119
rect 324 -120 325 -119
rect 325 -120 326 -119
rect 326 -120 327 -119
rect 327 -120 328 -119
rect 328 -120 329 -119
rect 329 -120 330 -119
rect 330 -120 331 -119
rect 331 -120 332 -119
rect 332 -120 333 -119
rect 333 -120 334 -119
rect 334 -120 335 -119
rect 335 -120 336 -119
rect 336 -120 337 -119
rect 337 -120 338 -119
rect 338 -120 339 -119
rect 339 -120 340 -119
rect 340 -120 341 -119
rect 341 -120 342 -119
rect 342 -120 343 -119
rect 343 -120 344 -119
rect 344 -120 345 -119
rect 345 -120 346 -119
rect 346 -120 347 -119
rect 347 -120 348 -119
rect 348 -120 349 -119
rect 349 -120 350 -119
rect 350 -120 351 -119
rect 351 -120 352 -119
rect 352 -120 353 -119
rect 353 -120 354 -119
rect 354 -120 355 -119
rect 355 -120 356 -119
rect 356 -120 357 -119
rect 357 -120 358 -119
rect 358 -120 359 -119
rect 359 -120 360 -119
rect 360 -120 361 -119
rect 361 -120 362 -119
rect 362 -120 363 -119
rect 363 -120 364 -119
rect 364 -120 365 -119
rect 365 -120 366 -119
rect 366 -120 367 -119
rect 367 -120 368 -119
rect 368 -120 369 -119
rect 369 -120 370 -119
rect 370 -120 371 -119
rect 371 -120 372 -119
rect 372 -120 373 -119
rect 373 -120 374 -119
rect 374 -120 375 -119
rect 375 -120 376 -119
rect 376 -120 377 -119
rect 377 -120 378 -119
rect 378 -120 379 -119
rect 379 -120 380 -119
rect 380 -120 381 -119
rect 381 -120 382 -119
rect 382 -120 383 -119
rect 383 -120 384 -119
rect 384 -120 385 -119
rect 385 -120 386 -119
rect 386 -120 387 -119
rect 387 -120 388 -119
rect 388 -120 389 -119
rect 389 -120 390 -119
rect 390 -120 391 -119
rect 391 -120 392 -119
rect 392 -120 393 -119
rect 393 -120 394 -119
rect 394 -120 395 -119
rect 395 -120 396 -119
rect 396 -120 397 -119
rect 397 -120 398 -119
rect 398 -120 399 -119
rect 399 -120 400 -119
rect 400 -120 401 -119
rect 401 -120 402 -119
rect 402 -120 403 -119
rect 403 -120 404 -119
rect 404 -120 405 -119
rect 405 -120 406 -119
rect 406 -120 407 -119
rect 407 -120 408 -119
rect 408 -120 409 -119
rect 409 -120 410 -119
rect 410 -120 411 -119
rect 411 -120 412 -119
rect 412 -120 413 -119
rect 413 -120 414 -119
rect 414 -120 415 -119
rect 415 -120 416 -119
rect 416 -120 417 -119
rect 417 -120 418 -119
rect 418 -120 419 -119
rect 419 -120 420 -119
rect 420 -120 421 -119
rect 421 -120 422 -119
rect 422 -120 423 -119
rect 423 -120 424 -119
rect 424 -120 425 -119
rect 425 -120 426 -119
rect 426 -120 427 -119
rect 427 -120 428 -119
rect 428 -120 429 -119
rect 429 -120 430 -119
rect 430 -120 431 -119
rect 431 -120 432 -119
rect 432 -120 433 -119
rect 433 -120 434 -119
rect 434 -120 435 -119
rect 435 -120 436 -119
rect 436 -120 437 -119
rect 437 -120 438 -119
rect 438 -120 439 -119
rect 439 -120 440 -119
rect 440 -120 441 -119
rect 441 -120 442 -119
rect 442 -120 443 -119
rect 443 -120 444 -119
rect 444 -120 445 -119
rect 445 -120 446 -119
rect 446 -120 447 -119
rect 447 -120 448 -119
rect 448 -120 449 -119
rect 449 -120 450 -119
rect 450 -120 451 -119
rect 451 -120 452 -119
rect 452 -120 453 -119
rect 453 -120 454 -119
rect 454 -120 455 -119
rect 455 -120 456 -119
rect 456 -120 457 -119
rect 457 -120 458 -119
rect 458 -120 459 -119
rect 459 -120 460 -119
rect 460 -120 461 -119
rect 461 -120 462 -119
rect 462 -120 463 -119
rect 463 -120 464 -119
rect 464 -120 465 -119
rect 465 -120 466 -119
rect 466 -120 467 -119
rect 467 -120 468 -119
rect 468 -120 469 -119
rect 469 -120 470 -119
rect 470 -120 471 -119
rect 471 -120 472 -119
rect 472 -120 473 -119
rect 473 -120 474 -119
rect 474 -120 475 -119
rect 475 -120 476 -119
rect 476 -120 477 -119
rect 477 -120 478 -119
rect 478 -120 479 -119
rect 479 -120 480 -119
rect 2 -121 3 -120
rect 3 -121 4 -120
rect 4 -121 5 -120
rect 5 -121 6 -120
rect 6 -121 7 -120
rect 7 -121 8 -120
rect 8 -121 9 -120
rect 24 -121 25 -120
rect 25 -121 26 -120
rect 26 -121 27 -120
rect 27 -121 28 -120
rect 28 -121 29 -120
rect 29 -121 30 -120
rect 30 -121 31 -120
rect 31 -121 32 -120
rect 32 -121 33 -120
rect 33 -121 34 -120
rect 34 -121 35 -120
rect 35 -121 36 -120
rect 36 -121 37 -120
rect 37 -121 38 -120
rect 38 -121 39 -120
rect 39 -121 40 -120
rect 40 -121 41 -120
rect 56 -121 57 -120
rect 57 -121 58 -120
rect 58 -121 59 -120
rect 59 -121 60 -120
rect 60 -121 61 -120
rect 61 -121 62 -120
rect 62 -121 63 -120
rect 63 -121 64 -120
rect 64 -121 65 -120
rect 65 -121 66 -120
rect 66 -121 67 -120
rect 67 -121 68 -120
rect 68 -121 69 -120
rect 69 -121 70 -120
rect 70 -121 71 -120
rect 71 -121 72 -120
rect 72 -121 73 -120
rect 88 -121 89 -120
rect 89 -121 90 -120
rect 90 -121 91 -120
rect 91 -121 92 -120
rect 92 -121 93 -120
rect 93 -121 94 -120
rect 94 -121 95 -120
rect 95 -121 96 -120
rect 96 -121 97 -120
rect 97 -121 98 -120
rect 98 -121 99 -120
rect 99 -121 100 -120
rect 100 -121 101 -120
rect 101 -121 102 -120
rect 102 -121 103 -120
rect 103 -121 104 -120
rect 104 -121 105 -120
rect 120 -121 121 -120
rect 121 -121 122 -120
rect 122 -121 123 -120
rect 123 -121 124 -120
rect 124 -121 125 -120
rect 125 -121 126 -120
rect 126 -121 127 -120
rect 127 -121 128 -120
rect 128 -121 129 -120
rect 129 -121 130 -120
rect 130 -121 131 -120
rect 131 -121 132 -120
rect 132 -121 133 -120
rect 133 -121 134 -120
rect 134 -121 135 -120
rect 135 -121 136 -120
rect 136 -121 137 -120
rect 152 -121 153 -120
rect 153 -121 154 -120
rect 154 -121 155 -120
rect 155 -121 156 -120
rect 156 -121 157 -120
rect 157 -121 158 -120
rect 158 -121 159 -120
rect 159 -121 160 -120
rect 160 -121 161 -120
rect 161 -121 162 -120
rect 162 -121 163 -120
rect 163 -121 164 -120
rect 164 -121 165 -120
rect 165 -121 166 -120
rect 166 -121 167 -120
rect 167 -121 168 -120
rect 168 -121 169 -120
rect 184 -121 185 -120
rect 185 -121 186 -120
rect 186 -121 187 -120
rect 187 -121 188 -120
rect 188 -121 189 -120
rect 189 -121 190 -120
rect 190 -121 191 -120
rect 191 -121 192 -120
rect 192 -121 193 -120
rect 193 -121 194 -120
rect 194 -121 195 -120
rect 195 -121 196 -120
rect 196 -121 197 -120
rect 197 -121 198 -120
rect 198 -121 199 -120
rect 199 -121 200 -120
rect 200 -121 201 -120
rect 201 -121 202 -120
rect 202 -121 203 -120
rect 203 -121 204 -120
rect 204 -121 205 -120
rect 205 -121 206 -120
rect 206 -121 207 -120
rect 207 -121 208 -120
rect 208 -121 209 -120
rect 209 -121 210 -120
rect 210 -121 211 -120
rect 211 -121 212 -120
rect 212 -121 213 -120
rect 213 -121 214 -120
rect 214 -121 215 -120
rect 215 -121 216 -120
rect 216 -121 217 -120
rect 217 -121 218 -120
rect 218 -121 219 -120
rect 219 -121 220 -120
rect 220 -121 221 -120
rect 221 -121 222 -120
rect 222 -121 223 -120
rect 223 -121 224 -120
rect 224 -121 225 -120
rect 225 -121 226 -120
rect 226 -121 227 -120
rect 227 -121 228 -120
rect 228 -121 229 -120
rect 229 -121 230 -120
rect 230 -121 231 -120
rect 231 -121 232 -120
rect 232 -121 233 -120
rect 233 -121 234 -120
rect 234 -121 235 -120
rect 235 -121 236 -120
rect 236 -121 237 -120
rect 237 -121 238 -120
rect 238 -121 239 -120
rect 239 -121 240 -120
rect 240 -121 241 -120
rect 241 -121 242 -120
rect 242 -121 243 -120
rect 243 -121 244 -120
rect 244 -121 245 -120
rect 245 -121 246 -120
rect 246 -121 247 -120
rect 247 -121 248 -120
rect 248 -121 249 -120
rect 249 -121 250 -120
rect 250 -121 251 -120
rect 251 -121 252 -120
rect 252 -121 253 -120
rect 253 -121 254 -120
rect 254 -121 255 -120
rect 255 -121 256 -120
rect 256 -121 257 -120
rect 257 -121 258 -120
rect 258 -121 259 -120
rect 259 -121 260 -120
rect 260 -121 261 -120
rect 261 -121 262 -120
rect 262 -121 263 -120
rect 263 -121 264 -120
rect 264 -121 265 -120
rect 265 -121 266 -120
rect 266 -121 267 -120
rect 267 -121 268 -120
rect 268 -121 269 -120
rect 269 -121 270 -120
rect 270 -121 271 -120
rect 271 -121 272 -120
rect 272 -121 273 -120
rect 273 -121 274 -120
rect 274 -121 275 -120
rect 275 -121 276 -120
rect 276 -121 277 -120
rect 277 -121 278 -120
rect 278 -121 279 -120
rect 279 -121 280 -120
rect 280 -121 281 -120
rect 281 -121 282 -120
rect 282 -121 283 -120
rect 283 -121 284 -120
rect 284 -121 285 -120
rect 285 -121 286 -120
rect 286 -121 287 -120
rect 287 -121 288 -120
rect 288 -121 289 -120
rect 289 -121 290 -120
rect 290 -121 291 -120
rect 291 -121 292 -120
rect 292 -121 293 -120
rect 293 -121 294 -120
rect 294 -121 295 -120
rect 295 -121 296 -120
rect 296 -121 297 -120
rect 297 -121 298 -120
rect 298 -121 299 -120
rect 299 -121 300 -120
rect 300 -121 301 -120
rect 301 -121 302 -120
rect 302 -121 303 -120
rect 303 -121 304 -120
rect 304 -121 305 -120
rect 305 -121 306 -120
rect 306 -121 307 -120
rect 307 -121 308 -120
rect 308 -121 309 -120
rect 309 -121 310 -120
rect 310 -121 311 -120
rect 311 -121 312 -120
rect 312 -121 313 -120
rect 313 -121 314 -120
rect 314 -121 315 -120
rect 315 -121 316 -120
rect 316 -121 317 -120
rect 317 -121 318 -120
rect 318 -121 319 -120
rect 319 -121 320 -120
rect 320 -121 321 -120
rect 321 -121 322 -120
rect 322 -121 323 -120
rect 323 -121 324 -120
rect 324 -121 325 -120
rect 325 -121 326 -120
rect 326 -121 327 -120
rect 327 -121 328 -120
rect 328 -121 329 -120
rect 329 -121 330 -120
rect 330 -121 331 -120
rect 331 -121 332 -120
rect 332 -121 333 -120
rect 333 -121 334 -120
rect 334 -121 335 -120
rect 335 -121 336 -120
rect 336 -121 337 -120
rect 337 -121 338 -120
rect 338 -121 339 -120
rect 339 -121 340 -120
rect 340 -121 341 -120
rect 341 -121 342 -120
rect 342 -121 343 -120
rect 343 -121 344 -120
rect 344 -121 345 -120
rect 345 -121 346 -120
rect 346 -121 347 -120
rect 347 -121 348 -120
rect 348 -121 349 -120
rect 349 -121 350 -120
rect 350 -121 351 -120
rect 351 -121 352 -120
rect 352 -121 353 -120
rect 353 -121 354 -120
rect 354 -121 355 -120
rect 355 -121 356 -120
rect 356 -121 357 -120
rect 357 -121 358 -120
rect 358 -121 359 -120
rect 359 -121 360 -120
rect 360 -121 361 -120
rect 361 -121 362 -120
rect 362 -121 363 -120
rect 363 -121 364 -120
rect 364 -121 365 -120
rect 365 -121 366 -120
rect 366 -121 367 -120
rect 367 -121 368 -120
rect 368 -121 369 -120
rect 369 -121 370 -120
rect 370 -121 371 -120
rect 371 -121 372 -120
rect 372 -121 373 -120
rect 373 -121 374 -120
rect 374 -121 375 -120
rect 375 -121 376 -120
rect 376 -121 377 -120
rect 377 -121 378 -120
rect 378 -121 379 -120
rect 379 -121 380 -120
rect 380 -121 381 -120
rect 381 -121 382 -120
rect 382 -121 383 -120
rect 383 -121 384 -120
rect 384 -121 385 -120
rect 385 -121 386 -120
rect 386 -121 387 -120
rect 387 -121 388 -120
rect 388 -121 389 -120
rect 389 -121 390 -120
rect 390 -121 391 -120
rect 391 -121 392 -120
rect 392 -121 393 -120
rect 393 -121 394 -120
rect 394 -121 395 -120
rect 395 -121 396 -120
rect 396 -121 397 -120
rect 397 -121 398 -120
rect 398 -121 399 -120
rect 399 -121 400 -120
rect 400 -121 401 -120
rect 401 -121 402 -120
rect 402 -121 403 -120
rect 403 -121 404 -120
rect 404 -121 405 -120
rect 405 -121 406 -120
rect 406 -121 407 -120
rect 407 -121 408 -120
rect 408 -121 409 -120
rect 409 -121 410 -120
rect 410 -121 411 -120
rect 411 -121 412 -120
rect 412 -121 413 -120
rect 413 -121 414 -120
rect 414 -121 415 -120
rect 415 -121 416 -120
rect 416 -121 417 -120
rect 417 -121 418 -120
rect 418 -121 419 -120
rect 419 -121 420 -120
rect 420 -121 421 -120
rect 421 -121 422 -120
rect 422 -121 423 -120
rect 423 -121 424 -120
rect 424 -121 425 -120
rect 425 -121 426 -120
rect 426 -121 427 -120
rect 427 -121 428 -120
rect 428 -121 429 -120
rect 429 -121 430 -120
rect 430 -121 431 -120
rect 431 -121 432 -120
rect 432 -121 433 -120
rect 433 -121 434 -120
rect 434 -121 435 -120
rect 435 -121 436 -120
rect 436 -121 437 -120
rect 437 -121 438 -120
rect 438 -121 439 -120
rect 439 -121 440 -120
rect 440 -121 441 -120
rect 441 -121 442 -120
rect 442 -121 443 -120
rect 443 -121 444 -120
rect 444 -121 445 -120
rect 445 -121 446 -120
rect 446 -121 447 -120
rect 447 -121 448 -120
rect 448 -121 449 -120
rect 449 -121 450 -120
rect 450 -121 451 -120
rect 451 -121 452 -120
rect 452 -121 453 -120
rect 453 -121 454 -120
rect 454 -121 455 -120
rect 455 -121 456 -120
rect 456 -121 457 -120
rect 457 -121 458 -120
rect 458 -121 459 -120
rect 459 -121 460 -120
rect 460 -121 461 -120
rect 461 -121 462 -120
rect 462 -121 463 -120
rect 463 -121 464 -120
rect 464 -121 465 -120
rect 465 -121 466 -120
rect 466 -121 467 -120
rect 467 -121 468 -120
rect 468 -121 469 -120
rect 469 -121 470 -120
rect 470 -121 471 -120
rect 471 -121 472 -120
rect 472 -121 473 -120
rect 473 -121 474 -120
rect 474 -121 475 -120
rect 475 -121 476 -120
rect 476 -121 477 -120
rect 477 -121 478 -120
rect 478 -121 479 -120
rect 479 -121 480 -120
rect 2 -122 3 -121
rect 3 -122 4 -121
rect 4 -122 5 -121
rect 5 -122 6 -121
rect 6 -122 7 -121
rect 7 -122 8 -121
rect 8 -122 9 -121
rect 9 -122 10 -121
rect 10 -122 11 -121
rect 23 -122 24 -121
rect 24 -122 25 -121
rect 25 -122 26 -121
rect 26 -122 27 -121
rect 27 -122 28 -121
rect 28 -122 29 -121
rect 29 -122 30 -121
rect 30 -122 31 -121
rect 31 -122 32 -121
rect 32 -122 33 -121
rect 33 -122 34 -121
rect 34 -122 35 -121
rect 35 -122 36 -121
rect 36 -122 37 -121
rect 37 -122 38 -121
rect 38 -122 39 -121
rect 39 -122 40 -121
rect 40 -122 41 -121
rect 41 -122 42 -121
rect 42 -122 43 -121
rect 55 -122 56 -121
rect 56 -122 57 -121
rect 57 -122 58 -121
rect 58 -122 59 -121
rect 59 -122 60 -121
rect 60 -122 61 -121
rect 61 -122 62 -121
rect 62 -122 63 -121
rect 63 -122 64 -121
rect 64 -122 65 -121
rect 65 -122 66 -121
rect 66 -122 67 -121
rect 67 -122 68 -121
rect 68 -122 69 -121
rect 69 -122 70 -121
rect 70 -122 71 -121
rect 71 -122 72 -121
rect 72 -122 73 -121
rect 73 -122 74 -121
rect 74 -122 75 -121
rect 87 -122 88 -121
rect 88 -122 89 -121
rect 89 -122 90 -121
rect 90 -122 91 -121
rect 91 -122 92 -121
rect 92 -122 93 -121
rect 93 -122 94 -121
rect 94 -122 95 -121
rect 95 -122 96 -121
rect 96 -122 97 -121
rect 97 -122 98 -121
rect 98 -122 99 -121
rect 99 -122 100 -121
rect 100 -122 101 -121
rect 101 -122 102 -121
rect 102 -122 103 -121
rect 103 -122 104 -121
rect 104 -122 105 -121
rect 105 -122 106 -121
rect 106 -122 107 -121
rect 119 -122 120 -121
rect 120 -122 121 -121
rect 121 -122 122 -121
rect 122 -122 123 -121
rect 123 -122 124 -121
rect 124 -122 125 -121
rect 125 -122 126 -121
rect 126 -122 127 -121
rect 127 -122 128 -121
rect 128 -122 129 -121
rect 129 -122 130 -121
rect 130 -122 131 -121
rect 131 -122 132 -121
rect 132 -122 133 -121
rect 133 -122 134 -121
rect 134 -122 135 -121
rect 135 -122 136 -121
rect 136 -122 137 -121
rect 137 -122 138 -121
rect 138 -122 139 -121
rect 151 -122 152 -121
rect 152 -122 153 -121
rect 153 -122 154 -121
rect 154 -122 155 -121
rect 155 -122 156 -121
rect 156 -122 157 -121
rect 157 -122 158 -121
rect 158 -122 159 -121
rect 159 -122 160 -121
rect 160 -122 161 -121
rect 161 -122 162 -121
rect 162 -122 163 -121
rect 163 -122 164 -121
rect 164 -122 165 -121
rect 165 -122 166 -121
rect 166 -122 167 -121
rect 167 -122 168 -121
rect 168 -122 169 -121
rect 169 -122 170 -121
rect 170 -122 171 -121
rect 183 -122 184 -121
rect 184 -122 185 -121
rect 185 -122 186 -121
rect 186 -122 187 -121
rect 187 -122 188 -121
rect 188 -122 189 -121
rect 189 -122 190 -121
rect 190 -122 191 -121
rect 191 -122 192 -121
rect 192 -122 193 -121
rect 193 -122 194 -121
rect 194 -122 195 -121
rect 195 -122 196 -121
rect 196 -122 197 -121
rect 197 -122 198 -121
rect 198 -122 199 -121
rect 199 -122 200 -121
rect 200 -122 201 -121
rect 201 -122 202 -121
rect 202 -122 203 -121
rect 203 -122 204 -121
rect 204 -122 205 -121
rect 205 -122 206 -121
rect 206 -122 207 -121
rect 207 -122 208 -121
rect 208 -122 209 -121
rect 209 -122 210 -121
rect 210 -122 211 -121
rect 211 -122 212 -121
rect 212 -122 213 -121
rect 213 -122 214 -121
rect 214 -122 215 -121
rect 215 -122 216 -121
rect 216 -122 217 -121
rect 217 -122 218 -121
rect 218 -122 219 -121
rect 219 -122 220 -121
rect 220 -122 221 -121
rect 221 -122 222 -121
rect 222 -122 223 -121
rect 223 -122 224 -121
rect 224 -122 225 -121
rect 225 -122 226 -121
rect 226 -122 227 -121
rect 227 -122 228 -121
rect 228 -122 229 -121
rect 229 -122 230 -121
rect 230 -122 231 -121
rect 231 -122 232 -121
rect 232 -122 233 -121
rect 233 -122 234 -121
rect 234 -122 235 -121
rect 235 -122 236 -121
rect 236 -122 237 -121
rect 237 -122 238 -121
rect 238 -122 239 -121
rect 239 -122 240 -121
rect 240 -122 241 -121
rect 241 -122 242 -121
rect 242 -122 243 -121
rect 243 -122 244 -121
rect 244 -122 245 -121
rect 245 -122 246 -121
rect 246 -122 247 -121
rect 247 -122 248 -121
rect 248 -122 249 -121
rect 249 -122 250 -121
rect 250 -122 251 -121
rect 251 -122 252 -121
rect 252 -122 253 -121
rect 253 -122 254 -121
rect 254 -122 255 -121
rect 255 -122 256 -121
rect 256 -122 257 -121
rect 257 -122 258 -121
rect 258 -122 259 -121
rect 259 -122 260 -121
rect 260 -122 261 -121
rect 261 -122 262 -121
rect 262 -122 263 -121
rect 263 -122 264 -121
rect 264 -122 265 -121
rect 265 -122 266 -121
rect 266 -122 267 -121
rect 267 -122 268 -121
rect 268 -122 269 -121
rect 269 -122 270 -121
rect 270 -122 271 -121
rect 271 -122 272 -121
rect 272 -122 273 -121
rect 273 -122 274 -121
rect 274 -122 275 -121
rect 275 -122 276 -121
rect 276 -122 277 -121
rect 277 -122 278 -121
rect 278 -122 279 -121
rect 279 -122 280 -121
rect 280 -122 281 -121
rect 281 -122 282 -121
rect 282 -122 283 -121
rect 283 -122 284 -121
rect 284 -122 285 -121
rect 285 -122 286 -121
rect 286 -122 287 -121
rect 287 -122 288 -121
rect 288 -122 289 -121
rect 289 -122 290 -121
rect 290 -122 291 -121
rect 291 -122 292 -121
rect 292 -122 293 -121
rect 293 -122 294 -121
rect 294 -122 295 -121
rect 295 -122 296 -121
rect 296 -122 297 -121
rect 297 -122 298 -121
rect 298 -122 299 -121
rect 299 -122 300 -121
rect 300 -122 301 -121
rect 301 -122 302 -121
rect 302 -122 303 -121
rect 303 -122 304 -121
rect 304 -122 305 -121
rect 305 -122 306 -121
rect 306 -122 307 -121
rect 307 -122 308 -121
rect 308 -122 309 -121
rect 309 -122 310 -121
rect 310 -122 311 -121
rect 311 -122 312 -121
rect 312 -122 313 -121
rect 313 -122 314 -121
rect 314 -122 315 -121
rect 315 -122 316 -121
rect 316 -122 317 -121
rect 317 -122 318 -121
rect 318 -122 319 -121
rect 319 -122 320 -121
rect 320 -122 321 -121
rect 321 -122 322 -121
rect 322 -122 323 -121
rect 323 -122 324 -121
rect 324 -122 325 -121
rect 325 -122 326 -121
rect 326 -122 327 -121
rect 327 -122 328 -121
rect 328 -122 329 -121
rect 329 -122 330 -121
rect 330 -122 331 -121
rect 331 -122 332 -121
rect 332 -122 333 -121
rect 333 -122 334 -121
rect 334 -122 335 -121
rect 335 -122 336 -121
rect 336 -122 337 -121
rect 337 -122 338 -121
rect 338 -122 339 -121
rect 339 -122 340 -121
rect 340 -122 341 -121
rect 341 -122 342 -121
rect 342 -122 343 -121
rect 343 -122 344 -121
rect 344 -122 345 -121
rect 345 -122 346 -121
rect 346 -122 347 -121
rect 347 -122 348 -121
rect 348 -122 349 -121
rect 349 -122 350 -121
rect 350 -122 351 -121
rect 351 -122 352 -121
rect 352 -122 353 -121
rect 353 -122 354 -121
rect 354 -122 355 -121
rect 355 -122 356 -121
rect 356 -122 357 -121
rect 357 -122 358 -121
rect 358 -122 359 -121
rect 359 -122 360 -121
rect 360 -122 361 -121
rect 361 -122 362 -121
rect 362 -122 363 -121
rect 363 -122 364 -121
rect 364 -122 365 -121
rect 365 -122 366 -121
rect 366 -122 367 -121
rect 367 -122 368 -121
rect 368 -122 369 -121
rect 369 -122 370 -121
rect 370 -122 371 -121
rect 371 -122 372 -121
rect 372 -122 373 -121
rect 373 -122 374 -121
rect 374 -122 375 -121
rect 375 -122 376 -121
rect 376 -122 377 -121
rect 377 -122 378 -121
rect 378 -122 379 -121
rect 379 -122 380 -121
rect 380 -122 381 -121
rect 381 -122 382 -121
rect 382 -122 383 -121
rect 383 -122 384 -121
rect 384 -122 385 -121
rect 385 -122 386 -121
rect 386 -122 387 -121
rect 387 -122 388 -121
rect 388 -122 389 -121
rect 389 -122 390 -121
rect 390 -122 391 -121
rect 391 -122 392 -121
rect 392 -122 393 -121
rect 393 -122 394 -121
rect 394 -122 395 -121
rect 395 -122 396 -121
rect 396 -122 397 -121
rect 397 -122 398 -121
rect 398 -122 399 -121
rect 399 -122 400 -121
rect 400 -122 401 -121
rect 401 -122 402 -121
rect 402 -122 403 -121
rect 403 -122 404 -121
rect 404 -122 405 -121
rect 405 -122 406 -121
rect 406 -122 407 -121
rect 407 -122 408 -121
rect 408 -122 409 -121
rect 409 -122 410 -121
rect 410 -122 411 -121
rect 411 -122 412 -121
rect 412 -122 413 -121
rect 413 -122 414 -121
rect 414 -122 415 -121
rect 415 -122 416 -121
rect 416 -122 417 -121
rect 417 -122 418 -121
rect 418 -122 419 -121
rect 419 -122 420 -121
rect 420 -122 421 -121
rect 421 -122 422 -121
rect 422 -122 423 -121
rect 423 -122 424 -121
rect 424 -122 425 -121
rect 425 -122 426 -121
rect 426 -122 427 -121
rect 427 -122 428 -121
rect 428 -122 429 -121
rect 429 -122 430 -121
rect 430 -122 431 -121
rect 431 -122 432 -121
rect 432 -122 433 -121
rect 433 -122 434 -121
rect 434 -122 435 -121
rect 435 -122 436 -121
rect 436 -122 437 -121
rect 437 -122 438 -121
rect 438 -122 439 -121
rect 439 -122 440 -121
rect 440 -122 441 -121
rect 441 -122 442 -121
rect 442 -122 443 -121
rect 443 -122 444 -121
rect 444 -122 445 -121
rect 445 -122 446 -121
rect 446 -122 447 -121
rect 447 -122 448 -121
rect 448 -122 449 -121
rect 449 -122 450 -121
rect 450 -122 451 -121
rect 451 -122 452 -121
rect 452 -122 453 -121
rect 453 -122 454 -121
rect 454 -122 455 -121
rect 455 -122 456 -121
rect 456 -122 457 -121
rect 457 -122 458 -121
rect 458 -122 459 -121
rect 459 -122 460 -121
rect 460 -122 461 -121
rect 461 -122 462 -121
rect 462 -122 463 -121
rect 463 -122 464 -121
rect 464 -122 465 -121
rect 465 -122 466 -121
rect 466 -122 467 -121
rect 467 -122 468 -121
rect 468 -122 469 -121
rect 469 -122 470 -121
rect 470 -122 471 -121
rect 471 -122 472 -121
rect 472 -122 473 -121
rect 473 -122 474 -121
rect 474 -122 475 -121
rect 475 -122 476 -121
rect 476 -122 477 -121
rect 477 -122 478 -121
rect 478 -122 479 -121
rect 479 -122 480 -121
rect 2 -123 3 -122
rect 3 -123 4 -122
rect 4 -123 5 -122
rect 5 -123 6 -122
rect 6 -123 7 -122
rect 7 -123 8 -122
rect 8 -123 9 -122
rect 9 -123 10 -122
rect 10 -123 11 -122
rect 11 -123 12 -122
rect 22 -123 23 -122
rect 23 -123 24 -122
rect 24 -123 25 -122
rect 25 -123 26 -122
rect 26 -123 27 -122
rect 27 -123 28 -122
rect 28 -123 29 -122
rect 29 -123 30 -122
rect 30 -123 31 -122
rect 31 -123 32 -122
rect 32 -123 33 -122
rect 33 -123 34 -122
rect 34 -123 35 -122
rect 35 -123 36 -122
rect 36 -123 37 -122
rect 37 -123 38 -122
rect 38 -123 39 -122
rect 39 -123 40 -122
rect 40 -123 41 -122
rect 41 -123 42 -122
rect 42 -123 43 -122
rect 43 -123 44 -122
rect 54 -123 55 -122
rect 55 -123 56 -122
rect 56 -123 57 -122
rect 57 -123 58 -122
rect 58 -123 59 -122
rect 59 -123 60 -122
rect 60 -123 61 -122
rect 61 -123 62 -122
rect 62 -123 63 -122
rect 63 -123 64 -122
rect 64 -123 65 -122
rect 65 -123 66 -122
rect 66 -123 67 -122
rect 67 -123 68 -122
rect 68 -123 69 -122
rect 69 -123 70 -122
rect 70 -123 71 -122
rect 71 -123 72 -122
rect 72 -123 73 -122
rect 73 -123 74 -122
rect 74 -123 75 -122
rect 75 -123 76 -122
rect 86 -123 87 -122
rect 87 -123 88 -122
rect 88 -123 89 -122
rect 89 -123 90 -122
rect 90 -123 91 -122
rect 91 -123 92 -122
rect 92 -123 93 -122
rect 93 -123 94 -122
rect 94 -123 95 -122
rect 95 -123 96 -122
rect 96 -123 97 -122
rect 97 -123 98 -122
rect 98 -123 99 -122
rect 99 -123 100 -122
rect 100 -123 101 -122
rect 101 -123 102 -122
rect 102 -123 103 -122
rect 103 -123 104 -122
rect 104 -123 105 -122
rect 105 -123 106 -122
rect 106 -123 107 -122
rect 107 -123 108 -122
rect 118 -123 119 -122
rect 119 -123 120 -122
rect 120 -123 121 -122
rect 121 -123 122 -122
rect 122 -123 123 -122
rect 123 -123 124 -122
rect 124 -123 125 -122
rect 125 -123 126 -122
rect 126 -123 127 -122
rect 127 -123 128 -122
rect 128 -123 129 -122
rect 129 -123 130 -122
rect 130 -123 131 -122
rect 131 -123 132 -122
rect 132 -123 133 -122
rect 133 -123 134 -122
rect 134 -123 135 -122
rect 135 -123 136 -122
rect 136 -123 137 -122
rect 137 -123 138 -122
rect 138 -123 139 -122
rect 139 -123 140 -122
rect 150 -123 151 -122
rect 151 -123 152 -122
rect 152 -123 153 -122
rect 153 -123 154 -122
rect 154 -123 155 -122
rect 155 -123 156 -122
rect 156 -123 157 -122
rect 157 -123 158 -122
rect 158 -123 159 -122
rect 159 -123 160 -122
rect 160 -123 161 -122
rect 161 -123 162 -122
rect 162 -123 163 -122
rect 163 -123 164 -122
rect 164 -123 165 -122
rect 165 -123 166 -122
rect 166 -123 167 -122
rect 167 -123 168 -122
rect 168 -123 169 -122
rect 169 -123 170 -122
rect 170 -123 171 -122
rect 171 -123 172 -122
rect 182 -123 183 -122
rect 183 -123 184 -122
rect 184 -123 185 -122
rect 185 -123 186 -122
rect 186 -123 187 -122
rect 187 -123 188 -122
rect 188 -123 189 -122
rect 189 -123 190 -122
rect 190 -123 191 -122
rect 191 -123 192 -122
rect 192 -123 193 -122
rect 193 -123 194 -122
rect 194 -123 195 -122
rect 195 -123 196 -122
rect 196 -123 197 -122
rect 197 -123 198 -122
rect 198 -123 199 -122
rect 199 -123 200 -122
rect 200 -123 201 -122
rect 201 -123 202 -122
rect 202 -123 203 -122
rect 203 -123 204 -122
rect 204 -123 205 -122
rect 205 -123 206 -122
rect 206 -123 207 -122
rect 207 -123 208 -122
rect 208 -123 209 -122
rect 209 -123 210 -122
rect 210 -123 211 -122
rect 211 -123 212 -122
rect 212 -123 213 -122
rect 213 -123 214 -122
rect 214 -123 215 -122
rect 215 -123 216 -122
rect 216 -123 217 -122
rect 217 -123 218 -122
rect 218 -123 219 -122
rect 219 -123 220 -122
rect 220 -123 221 -122
rect 221 -123 222 -122
rect 222 -123 223 -122
rect 223 -123 224 -122
rect 224 -123 225 -122
rect 225 -123 226 -122
rect 226 -123 227 -122
rect 227 -123 228 -122
rect 228 -123 229 -122
rect 229 -123 230 -122
rect 230 -123 231 -122
rect 231 -123 232 -122
rect 232 -123 233 -122
rect 233 -123 234 -122
rect 234 -123 235 -122
rect 235 -123 236 -122
rect 236 -123 237 -122
rect 237 -123 238 -122
rect 238 -123 239 -122
rect 239 -123 240 -122
rect 240 -123 241 -122
rect 241 -123 242 -122
rect 242 -123 243 -122
rect 243 -123 244 -122
rect 244 -123 245 -122
rect 245 -123 246 -122
rect 246 -123 247 -122
rect 247 -123 248 -122
rect 248 -123 249 -122
rect 249 -123 250 -122
rect 250 -123 251 -122
rect 251 -123 252 -122
rect 252 -123 253 -122
rect 253 -123 254 -122
rect 254 -123 255 -122
rect 255 -123 256 -122
rect 256 -123 257 -122
rect 257 -123 258 -122
rect 258 -123 259 -122
rect 259 -123 260 -122
rect 260 -123 261 -122
rect 261 -123 262 -122
rect 262 -123 263 -122
rect 263 -123 264 -122
rect 264 -123 265 -122
rect 265 -123 266 -122
rect 266 -123 267 -122
rect 267 -123 268 -122
rect 268 -123 269 -122
rect 269 -123 270 -122
rect 270 -123 271 -122
rect 271 -123 272 -122
rect 272 -123 273 -122
rect 273 -123 274 -122
rect 274 -123 275 -122
rect 275 -123 276 -122
rect 276 -123 277 -122
rect 277 -123 278 -122
rect 278 -123 279 -122
rect 279 -123 280 -122
rect 280 -123 281 -122
rect 281 -123 282 -122
rect 282 -123 283 -122
rect 283 -123 284 -122
rect 284 -123 285 -122
rect 285 -123 286 -122
rect 286 -123 287 -122
rect 287 -123 288 -122
rect 288 -123 289 -122
rect 289 -123 290 -122
rect 290 -123 291 -122
rect 291 -123 292 -122
rect 292 -123 293 -122
rect 293 -123 294 -122
rect 294 -123 295 -122
rect 295 -123 296 -122
rect 296 -123 297 -122
rect 297 -123 298 -122
rect 298 -123 299 -122
rect 299 -123 300 -122
rect 300 -123 301 -122
rect 301 -123 302 -122
rect 302 -123 303 -122
rect 303 -123 304 -122
rect 304 -123 305 -122
rect 305 -123 306 -122
rect 306 -123 307 -122
rect 307 -123 308 -122
rect 308 -123 309 -122
rect 309 -123 310 -122
rect 310 -123 311 -122
rect 311 -123 312 -122
rect 312 -123 313 -122
rect 313 -123 314 -122
rect 314 -123 315 -122
rect 315 -123 316 -122
rect 316 -123 317 -122
rect 317 -123 318 -122
rect 318 -123 319 -122
rect 319 -123 320 -122
rect 320 -123 321 -122
rect 321 -123 322 -122
rect 322 -123 323 -122
rect 323 -123 324 -122
rect 324 -123 325 -122
rect 325 -123 326 -122
rect 326 -123 327 -122
rect 327 -123 328 -122
rect 328 -123 329 -122
rect 329 -123 330 -122
rect 330 -123 331 -122
rect 331 -123 332 -122
rect 332 -123 333 -122
rect 333 -123 334 -122
rect 334 -123 335 -122
rect 335 -123 336 -122
rect 336 -123 337 -122
rect 337 -123 338 -122
rect 338 -123 339 -122
rect 339 -123 340 -122
rect 340 -123 341 -122
rect 341 -123 342 -122
rect 342 -123 343 -122
rect 343 -123 344 -122
rect 344 -123 345 -122
rect 345 -123 346 -122
rect 346 -123 347 -122
rect 347 -123 348 -122
rect 348 -123 349 -122
rect 349 -123 350 -122
rect 350 -123 351 -122
rect 351 -123 352 -122
rect 352 -123 353 -122
rect 353 -123 354 -122
rect 354 -123 355 -122
rect 355 -123 356 -122
rect 356 -123 357 -122
rect 357 -123 358 -122
rect 358 -123 359 -122
rect 359 -123 360 -122
rect 360 -123 361 -122
rect 361 -123 362 -122
rect 362 -123 363 -122
rect 363 -123 364 -122
rect 364 -123 365 -122
rect 365 -123 366 -122
rect 366 -123 367 -122
rect 367 -123 368 -122
rect 368 -123 369 -122
rect 369 -123 370 -122
rect 370 -123 371 -122
rect 371 -123 372 -122
rect 372 -123 373 -122
rect 373 -123 374 -122
rect 374 -123 375 -122
rect 375 -123 376 -122
rect 376 -123 377 -122
rect 377 -123 378 -122
rect 378 -123 379 -122
rect 379 -123 380 -122
rect 380 -123 381 -122
rect 381 -123 382 -122
rect 382 -123 383 -122
rect 383 -123 384 -122
rect 384 -123 385 -122
rect 385 -123 386 -122
rect 386 -123 387 -122
rect 387 -123 388 -122
rect 388 -123 389 -122
rect 389 -123 390 -122
rect 390 -123 391 -122
rect 391 -123 392 -122
rect 392 -123 393 -122
rect 393 -123 394 -122
rect 394 -123 395 -122
rect 395 -123 396 -122
rect 396 -123 397 -122
rect 397 -123 398 -122
rect 398 -123 399 -122
rect 399 -123 400 -122
rect 400 -123 401 -122
rect 401 -123 402 -122
rect 402 -123 403 -122
rect 403 -123 404 -122
rect 404 -123 405 -122
rect 405 -123 406 -122
rect 406 -123 407 -122
rect 407 -123 408 -122
rect 408 -123 409 -122
rect 409 -123 410 -122
rect 410 -123 411 -122
rect 411 -123 412 -122
rect 412 -123 413 -122
rect 413 -123 414 -122
rect 414 -123 415 -122
rect 415 -123 416 -122
rect 416 -123 417 -122
rect 417 -123 418 -122
rect 418 -123 419 -122
rect 419 -123 420 -122
rect 420 -123 421 -122
rect 421 -123 422 -122
rect 422 -123 423 -122
rect 423 -123 424 -122
rect 424 -123 425 -122
rect 425 -123 426 -122
rect 426 -123 427 -122
rect 427 -123 428 -122
rect 428 -123 429 -122
rect 429 -123 430 -122
rect 430 -123 431 -122
rect 431 -123 432 -122
rect 432 -123 433 -122
rect 433 -123 434 -122
rect 434 -123 435 -122
rect 435 -123 436 -122
rect 436 -123 437 -122
rect 437 -123 438 -122
rect 438 -123 439 -122
rect 439 -123 440 -122
rect 440 -123 441 -122
rect 441 -123 442 -122
rect 442 -123 443 -122
rect 443 -123 444 -122
rect 444 -123 445 -122
rect 445 -123 446 -122
rect 446 -123 447 -122
rect 447 -123 448 -122
rect 448 -123 449 -122
rect 449 -123 450 -122
rect 450 -123 451 -122
rect 451 -123 452 -122
rect 452 -123 453 -122
rect 453 -123 454 -122
rect 454 -123 455 -122
rect 455 -123 456 -122
rect 456 -123 457 -122
rect 457 -123 458 -122
rect 458 -123 459 -122
rect 459 -123 460 -122
rect 460 -123 461 -122
rect 461 -123 462 -122
rect 462 -123 463 -122
rect 463 -123 464 -122
rect 464 -123 465 -122
rect 465 -123 466 -122
rect 466 -123 467 -122
rect 467 -123 468 -122
rect 468 -123 469 -122
rect 469 -123 470 -122
rect 470 -123 471 -122
rect 471 -123 472 -122
rect 472 -123 473 -122
rect 473 -123 474 -122
rect 474 -123 475 -122
rect 475 -123 476 -122
rect 476 -123 477 -122
rect 477 -123 478 -122
rect 478 -123 479 -122
rect 479 -123 480 -122
rect 2 -124 3 -123
rect 3 -124 4 -123
rect 4 -124 5 -123
rect 5 -124 6 -123
rect 6 -124 7 -123
rect 7 -124 8 -123
rect 8 -124 9 -123
rect 9 -124 10 -123
rect 10 -124 11 -123
rect 11 -124 12 -123
rect 21 -124 22 -123
rect 22 -124 23 -123
rect 23 -124 24 -123
rect 24 -124 25 -123
rect 25 -124 26 -123
rect 26 -124 27 -123
rect 27 -124 28 -123
rect 28 -124 29 -123
rect 29 -124 30 -123
rect 30 -124 31 -123
rect 31 -124 32 -123
rect 32 -124 33 -123
rect 33 -124 34 -123
rect 34 -124 35 -123
rect 35 -124 36 -123
rect 36 -124 37 -123
rect 37 -124 38 -123
rect 38 -124 39 -123
rect 39 -124 40 -123
rect 40 -124 41 -123
rect 41 -124 42 -123
rect 42 -124 43 -123
rect 43 -124 44 -123
rect 53 -124 54 -123
rect 54 -124 55 -123
rect 55 -124 56 -123
rect 56 -124 57 -123
rect 57 -124 58 -123
rect 58 -124 59 -123
rect 59 -124 60 -123
rect 60 -124 61 -123
rect 61 -124 62 -123
rect 62 -124 63 -123
rect 63 -124 64 -123
rect 64 -124 65 -123
rect 65 -124 66 -123
rect 66 -124 67 -123
rect 67 -124 68 -123
rect 68 -124 69 -123
rect 69 -124 70 -123
rect 70 -124 71 -123
rect 71 -124 72 -123
rect 72 -124 73 -123
rect 73 -124 74 -123
rect 74 -124 75 -123
rect 75 -124 76 -123
rect 85 -124 86 -123
rect 86 -124 87 -123
rect 87 -124 88 -123
rect 88 -124 89 -123
rect 89 -124 90 -123
rect 90 -124 91 -123
rect 91 -124 92 -123
rect 92 -124 93 -123
rect 93 -124 94 -123
rect 94 -124 95 -123
rect 95 -124 96 -123
rect 96 -124 97 -123
rect 97 -124 98 -123
rect 98 -124 99 -123
rect 99 -124 100 -123
rect 100 -124 101 -123
rect 101 -124 102 -123
rect 102 -124 103 -123
rect 103 -124 104 -123
rect 104 -124 105 -123
rect 105 -124 106 -123
rect 106 -124 107 -123
rect 107 -124 108 -123
rect 117 -124 118 -123
rect 118 -124 119 -123
rect 119 -124 120 -123
rect 120 -124 121 -123
rect 121 -124 122 -123
rect 122 -124 123 -123
rect 123 -124 124 -123
rect 124 -124 125 -123
rect 125 -124 126 -123
rect 126 -124 127 -123
rect 127 -124 128 -123
rect 128 -124 129 -123
rect 129 -124 130 -123
rect 130 -124 131 -123
rect 131 -124 132 -123
rect 132 -124 133 -123
rect 133 -124 134 -123
rect 134 -124 135 -123
rect 135 -124 136 -123
rect 136 -124 137 -123
rect 137 -124 138 -123
rect 138 -124 139 -123
rect 139 -124 140 -123
rect 149 -124 150 -123
rect 150 -124 151 -123
rect 151 -124 152 -123
rect 152 -124 153 -123
rect 153 -124 154 -123
rect 154 -124 155 -123
rect 155 -124 156 -123
rect 156 -124 157 -123
rect 157 -124 158 -123
rect 158 -124 159 -123
rect 159 -124 160 -123
rect 160 -124 161 -123
rect 161 -124 162 -123
rect 162 -124 163 -123
rect 163 -124 164 -123
rect 164 -124 165 -123
rect 165 -124 166 -123
rect 166 -124 167 -123
rect 167 -124 168 -123
rect 168 -124 169 -123
rect 169 -124 170 -123
rect 170 -124 171 -123
rect 171 -124 172 -123
rect 181 -124 182 -123
rect 182 -124 183 -123
rect 183 -124 184 -123
rect 184 -124 185 -123
rect 185 -124 186 -123
rect 186 -124 187 -123
rect 187 -124 188 -123
rect 188 -124 189 -123
rect 189 -124 190 -123
rect 190 -124 191 -123
rect 191 -124 192 -123
rect 192 -124 193 -123
rect 193 -124 194 -123
rect 194 -124 195 -123
rect 195 -124 196 -123
rect 196 -124 197 -123
rect 197 -124 198 -123
rect 198 -124 199 -123
rect 199 -124 200 -123
rect 200 -124 201 -123
rect 201 -124 202 -123
rect 202 -124 203 -123
rect 203 -124 204 -123
rect 204 -124 205 -123
rect 205 -124 206 -123
rect 206 -124 207 -123
rect 207 -124 208 -123
rect 208 -124 209 -123
rect 209 -124 210 -123
rect 210 -124 211 -123
rect 211 -124 212 -123
rect 212 -124 213 -123
rect 213 -124 214 -123
rect 214 -124 215 -123
rect 215 -124 216 -123
rect 216 -124 217 -123
rect 217 -124 218 -123
rect 218 -124 219 -123
rect 219 -124 220 -123
rect 220 -124 221 -123
rect 221 -124 222 -123
rect 222 -124 223 -123
rect 223 -124 224 -123
rect 224 -124 225 -123
rect 225 -124 226 -123
rect 226 -124 227 -123
rect 227 -124 228 -123
rect 228 -124 229 -123
rect 229 -124 230 -123
rect 230 -124 231 -123
rect 231 -124 232 -123
rect 232 -124 233 -123
rect 233 -124 234 -123
rect 234 -124 235 -123
rect 235 -124 236 -123
rect 236 -124 237 -123
rect 237 -124 238 -123
rect 238 -124 239 -123
rect 239 -124 240 -123
rect 240 -124 241 -123
rect 241 -124 242 -123
rect 242 -124 243 -123
rect 243 -124 244 -123
rect 244 -124 245 -123
rect 245 -124 246 -123
rect 246 -124 247 -123
rect 247 -124 248 -123
rect 248 -124 249 -123
rect 249 -124 250 -123
rect 250 -124 251 -123
rect 251 -124 252 -123
rect 252 -124 253 -123
rect 253 -124 254 -123
rect 254 -124 255 -123
rect 255 -124 256 -123
rect 256 -124 257 -123
rect 257 -124 258 -123
rect 258 -124 259 -123
rect 259 -124 260 -123
rect 260 -124 261 -123
rect 261 -124 262 -123
rect 262 -124 263 -123
rect 263 -124 264 -123
rect 264 -124 265 -123
rect 265 -124 266 -123
rect 266 -124 267 -123
rect 267 -124 268 -123
rect 268 -124 269 -123
rect 269 -124 270 -123
rect 270 -124 271 -123
rect 271 -124 272 -123
rect 272 -124 273 -123
rect 273 -124 274 -123
rect 274 -124 275 -123
rect 275 -124 276 -123
rect 276 -124 277 -123
rect 277 -124 278 -123
rect 278 -124 279 -123
rect 279 -124 280 -123
rect 280 -124 281 -123
rect 281 -124 282 -123
rect 282 -124 283 -123
rect 283 -124 284 -123
rect 284 -124 285 -123
rect 285 -124 286 -123
rect 286 -124 287 -123
rect 287 -124 288 -123
rect 288 -124 289 -123
rect 289 -124 290 -123
rect 290 -124 291 -123
rect 291 -124 292 -123
rect 292 -124 293 -123
rect 293 -124 294 -123
rect 294 -124 295 -123
rect 295 -124 296 -123
rect 296 -124 297 -123
rect 297 -124 298 -123
rect 298 -124 299 -123
rect 299 -124 300 -123
rect 300 -124 301 -123
rect 301 -124 302 -123
rect 302 -124 303 -123
rect 303 -124 304 -123
rect 304 -124 305 -123
rect 305 -124 306 -123
rect 306 -124 307 -123
rect 307 -124 308 -123
rect 308 -124 309 -123
rect 309 -124 310 -123
rect 310 -124 311 -123
rect 311 -124 312 -123
rect 312 -124 313 -123
rect 313 -124 314 -123
rect 314 -124 315 -123
rect 315 -124 316 -123
rect 316 -124 317 -123
rect 317 -124 318 -123
rect 318 -124 319 -123
rect 319 -124 320 -123
rect 320 -124 321 -123
rect 321 -124 322 -123
rect 322 -124 323 -123
rect 323 -124 324 -123
rect 324 -124 325 -123
rect 325 -124 326 -123
rect 326 -124 327 -123
rect 327 -124 328 -123
rect 328 -124 329 -123
rect 329 -124 330 -123
rect 330 -124 331 -123
rect 331 -124 332 -123
rect 332 -124 333 -123
rect 333 -124 334 -123
rect 334 -124 335 -123
rect 335 -124 336 -123
rect 336 -124 337 -123
rect 337 -124 338 -123
rect 338 -124 339 -123
rect 339 -124 340 -123
rect 340 -124 341 -123
rect 341 -124 342 -123
rect 342 -124 343 -123
rect 343 -124 344 -123
rect 344 -124 345 -123
rect 345 -124 346 -123
rect 346 -124 347 -123
rect 347 -124 348 -123
rect 348 -124 349 -123
rect 349 -124 350 -123
rect 350 -124 351 -123
rect 351 -124 352 -123
rect 352 -124 353 -123
rect 353 -124 354 -123
rect 354 -124 355 -123
rect 355 -124 356 -123
rect 356 -124 357 -123
rect 357 -124 358 -123
rect 358 -124 359 -123
rect 359 -124 360 -123
rect 360 -124 361 -123
rect 361 -124 362 -123
rect 362 -124 363 -123
rect 363 -124 364 -123
rect 364 -124 365 -123
rect 365 -124 366 -123
rect 366 -124 367 -123
rect 367 -124 368 -123
rect 368 -124 369 -123
rect 369 -124 370 -123
rect 370 -124 371 -123
rect 371 -124 372 -123
rect 372 -124 373 -123
rect 373 -124 374 -123
rect 374 -124 375 -123
rect 375 -124 376 -123
rect 376 -124 377 -123
rect 377 -124 378 -123
rect 378 -124 379 -123
rect 379 -124 380 -123
rect 380 -124 381 -123
rect 381 -124 382 -123
rect 382 -124 383 -123
rect 383 -124 384 -123
rect 384 -124 385 -123
rect 385 -124 386 -123
rect 386 -124 387 -123
rect 387 -124 388 -123
rect 388 -124 389 -123
rect 389 -124 390 -123
rect 390 -124 391 -123
rect 391 -124 392 -123
rect 392 -124 393 -123
rect 393 -124 394 -123
rect 394 -124 395 -123
rect 395 -124 396 -123
rect 396 -124 397 -123
rect 397 -124 398 -123
rect 398 -124 399 -123
rect 399 -124 400 -123
rect 400 -124 401 -123
rect 401 -124 402 -123
rect 402 -124 403 -123
rect 403 -124 404 -123
rect 404 -124 405 -123
rect 405 -124 406 -123
rect 406 -124 407 -123
rect 407 -124 408 -123
rect 408 -124 409 -123
rect 409 -124 410 -123
rect 410 -124 411 -123
rect 411 -124 412 -123
rect 412 -124 413 -123
rect 413 -124 414 -123
rect 414 -124 415 -123
rect 415 -124 416 -123
rect 416 -124 417 -123
rect 417 -124 418 -123
rect 418 -124 419 -123
rect 419 -124 420 -123
rect 420 -124 421 -123
rect 421 -124 422 -123
rect 422 -124 423 -123
rect 423 -124 424 -123
rect 424 -124 425 -123
rect 425 -124 426 -123
rect 426 -124 427 -123
rect 427 -124 428 -123
rect 428 -124 429 -123
rect 429 -124 430 -123
rect 430 -124 431 -123
rect 431 -124 432 -123
rect 432 -124 433 -123
rect 433 -124 434 -123
rect 434 -124 435 -123
rect 435 -124 436 -123
rect 436 -124 437 -123
rect 437 -124 438 -123
rect 438 -124 439 -123
rect 439 -124 440 -123
rect 440 -124 441 -123
rect 441 -124 442 -123
rect 442 -124 443 -123
rect 443 -124 444 -123
rect 444 -124 445 -123
rect 445 -124 446 -123
rect 446 -124 447 -123
rect 447 -124 448 -123
rect 448 -124 449 -123
rect 449 -124 450 -123
rect 450 -124 451 -123
rect 451 -124 452 -123
rect 452 -124 453 -123
rect 453 -124 454 -123
rect 454 -124 455 -123
rect 455 -124 456 -123
rect 456 -124 457 -123
rect 457 -124 458 -123
rect 458 -124 459 -123
rect 459 -124 460 -123
rect 460 -124 461 -123
rect 461 -124 462 -123
rect 462 -124 463 -123
rect 463 -124 464 -123
rect 464 -124 465 -123
rect 465 -124 466 -123
rect 466 -124 467 -123
rect 467 -124 468 -123
rect 468 -124 469 -123
rect 469 -124 470 -123
rect 470 -124 471 -123
rect 471 -124 472 -123
rect 472 -124 473 -123
rect 473 -124 474 -123
rect 474 -124 475 -123
rect 475 -124 476 -123
rect 476 -124 477 -123
rect 477 -124 478 -123
rect 478 -124 479 -123
rect 479 -124 480 -123
rect 2 -125 3 -124
rect 3 -125 4 -124
rect 4 -125 5 -124
rect 5 -125 6 -124
rect 6 -125 7 -124
rect 7 -125 8 -124
rect 8 -125 9 -124
rect 9 -125 10 -124
rect 10 -125 11 -124
rect 11 -125 12 -124
rect 21 -125 22 -124
rect 22 -125 23 -124
rect 23 -125 24 -124
rect 24 -125 25 -124
rect 25 -125 26 -124
rect 26 -125 27 -124
rect 27 -125 28 -124
rect 28 -125 29 -124
rect 29 -125 30 -124
rect 30 -125 31 -124
rect 31 -125 32 -124
rect 32 -125 33 -124
rect 33 -125 34 -124
rect 34 -125 35 -124
rect 35 -125 36 -124
rect 36 -125 37 -124
rect 37 -125 38 -124
rect 38 -125 39 -124
rect 39 -125 40 -124
rect 40 -125 41 -124
rect 41 -125 42 -124
rect 42 -125 43 -124
rect 43 -125 44 -124
rect 53 -125 54 -124
rect 54 -125 55 -124
rect 55 -125 56 -124
rect 56 -125 57 -124
rect 57 -125 58 -124
rect 58 -125 59 -124
rect 59 -125 60 -124
rect 60 -125 61 -124
rect 61 -125 62 -124
rect 62 -125 63 -124
rect 63 -125 64 -124
rect 64 -125 65 -124
rect 65 -125 66 -124
rect 66 -125 67 -124
rect 67 -125 68 -124
rect 68 -125 69 -124
rect 69 -125 70 -124
rect 70 -125 71 -124
rect 71 -125 72 -124
rect 72 -125 73 -124
rect 73 -125 74 -124
rect 74 -125 75 -124
rect 75 -125 76 -124
rect 85 -125 86 -124
rect 86 -125 87 -124
rect 87 -125 88 -124
rect 88 -125 89 -124
rect 89 -125 90 -124
rect 90 -125 91 -124
rect 91 -125 92 -124
rect 92 -125 93 -124
rect 93 -125 94 -124
rect 94 -125 95 -124
rect 95 -125 96 -124
rect 96 -125 97 -124
rect 97 -125 98 -124
rect 98 -125 99 -124
rect 99 -125 100 -124
rect 100 -125 101 -124
rect 101 -125 102 -124
rect 102 -125 103 -124
rect 103 -125 104 -124
rect 104 -125 105 -124
rect 105 -125 106 -124
rect 106 -125 107 -124
rect 107 -125 108 -124
rect 117 -125 118 -124
rect 118 -125 119 -124
rect 119 -125 120 -124
rect 120 -125 121 -124
rect 121 -125 122 -124
rect 122 -125 123 -124
rect 123 -125 124 -124
rect 124 -125 125 -124
rect 125 -125 126 -124
rect 126 -125 127 -124
rect 127 -125 128 -124
rect 128 -125 129 -124
rect 129 -125 130 -124
rect 130 -125 131 -124
rect 131 -125 132 -124
rect 132 -125 133 -124
rect 133 -125 134 -124
rect 134 -125 135 -124
rect 135 -125 136 -124
rect 136 -125 137 -124
rect 137 -125 138 -124
rect 138 -125 139 -124
rect 139 -125 140 -124
rect 149 -125 150 -124
rect 150 -125 151 -124
rect 151 -125 152 -124
rect 152 -125 153 -124
rect 153 -125 154 -124
rect 154 -125 155 -124
rect 155 -125 156 -124
rect 156 -125 157 -124
rect 157 -125 158 -124
rect 158 -125 159 -124
rect 159 -125 160 -124
rect 160 -125 161 -124
rect 161 -125 162 -124
rect 162 -125 163 -124
rect 163 -125 164 -124
rect 164 -125 165 -124
rect 165 -125 166 -124
rect 166 -125 167 -124
rect 167 -125 168 -124
rect 168 -125 169 -124
rect 169 -125 170 -124
rect 170 -125 171 -124
rect 171 -125 172 -124
rect 181 -125 182 -124
rect 182 -125 183 -124
rect 183 -125 184 -124
rect 184 -125 185 -124
rect 185 -125 186 -124
rect 186 -125 187 -124
rect 187 -125 188 -124
rect 188 -125 189 -124
rect 189 -125 190 -124
rect 190 -125 191 -124
rect 191 -125 192 -124
rect 192 -125 193 -124
rect 193 -125 194 -124
rect 194 -125 195 -124
rect 195 -125 196 -124
rect 196 -125 197 -124
rect 197 -125 198 -124
rect 198 -125 199 -124
rect 199 -125 200 -124
rect 200 -125 201 -124
rect 201 -125 202 -124
rect 202 -125 203 -124
rect 203 -125 204 -124
rect 204 -125 205 -124
rect 205 -125 206 -124
rect 206 -125 207 -124
rect 207 -125 208 -124
rect 208 -125 209 -124
rect 209 -125 210 -124
rect 210 -125 211 -124
rect 211 -125 212 -124
rect 212 -125 213 -124
rect 213 -125 214 -124
rect 214 -125 215 -124
rect 215 -125 216 -124
rect 216 -125 217 -124
rect 217 -125 218 -124
rect 218 -125 219 -124
rect 219 -125 220 -124
rect 220 -125 221 -124
rect 221 -125 222 -124
rect 222 -125 223 -124
rect 223 -125 224 -124
rect 224 -125 225 -124
rect 225 -125 226 -124
rect 226 -125 227 -124
rect 227 -125 228 -124
rect 228 -125 229 -124
rect 229 -125 230 -124
rect 230 -125 231 -124
rect 231 -125 232 -124
rect 232 -125 233 -124
rect 233 -125 234 -124
rect 234 -125 235 -124
rect 235 -125 236 -124
rect 236 -125 237 -124
rect 237 -125 238 -124
rect 238 -125 239 -124
rect 239 -125 240 -124
rect 240 -125 241 -124
rect 241 -125 242 -124
rect 242 -125 243 -124
rect 243 -125 244 -124
rect 244 -125 245 -124
rect 245 -125 246 -124
rect 246 -125 247 -124
rect 247 -125 248 -124
rect 248 -125 249 -124
rect 249 -125 250 -124
rect 250 -125 251 -124
rect 251 -125 252 -124
rect 252 -125 253 -124
rect 253 -125 254 -124
rect 254 -125 255 -124
rect 255 -125 256 -124
rect 256 -125 257 -124
rect 257 -125 258 -124
rect 258 -125 259 -124
rect 259 -125 260 -124
rect 260 -125 261 -124
rect 261 -125 262 -124
rect 262 -125 263 -124
rect 263 -125 264 -124
rect 264 -125 265 -124
rect 265 -125 266 -124
rect 266 -125 267 -124
rect 267 -125 268 -124
rect 268 -125 269 -124
rect 269 -125 270 -124
rect 270 -125 271 -124
rect 271 -125 272 -124
rect 272 -125 273 -124
rect 273 -125 274 -124
rect 274 -125 275 -124
rect 275 -125 276 -124
rect 276 -125 277 -124
rect 277 -125 278 -124
rect 278 -125 279 -124
rect 279 -125 280 -124
rect 280 -125 281 -124
rect 281 -125 282 -124
rect 282 -125 283 -124
rect 283 -125 284 -124
rect 284 -125 285 -124
rect 285 -125 286 -124
rect 286 -125 287 -124
rect 287 -125 288 -124
rect 288 -125 289 -124
rect 289 -125 290 -124
rect 290 -125 291 -124
rect 291 -125 292 -124
rect 292 -125 293 -124
rect 293 -125 294 -124
rect 294 -125 295 -124
rect 295 -125 296 -124
rect 296 -125 297 -124
rect 297 -125 298 -124
rect 298 -125 299 -124
rect 299 -125 300 -124
rect 300 -125 301 -124
rect 301 -125 302 -124
rect 302 -125 303 -124
rect 303 -125 304 -124
rect 304 -125 305 -124
rect 305 -125 306 -124
rect 306 -125 307 -124
rect 307 -125 308 -124
rect 308 -125 309 -124
rect 309 -125 310 -124
rect 310 -125 311 -124
rect 311 -125 312 -124
rect 312 -125 313 -124
rect 313 -125 314 -124
rect 314 -125 315 -124
rect 315 -125 316 -124
rect 316 -125 317 -124
rect 317 -125 318 -124
rect 318 -125 319 -124
rect 319 -125 320 -124
rect 320 -125 321 -124
rect 321 -125 322 -124
rect 322 -125 323 -124
rect 323 -125 324 -124
rect 324 -125 325 -124
rect 325 -125 326 -124
rect 326 -125 327 -124
rect 327 -125 328 -124
rect 328 -125 329 -124
rect 329 -125 330 -124
rect 330 -125 331 -124
rect 331 -125 332 -124
rect 332 -125 333 -124
rect 333 -125 334 -124
rect 334 -125 335 -124
rect 335 -125 336 -124
rect 336 -125 337 -124
rect 337 -125 338 -124
rect 338 -125 339 -124
rect 339 -125 340 -124
rect 340 -125 341 -124
rect 341 -125 342 -124
rect 342 -125 343 -124
rect 343 -125 344 -124
rect 344 -125 345 -124
rect 345 -125 346 -124
rect 346 -125 347 -124
rect 347 -125 348 -124
rect 348 -125 349 -124
rect 349 -125 350 -124
rect 350 -125 351 -124
rect 351 -125 352 -124
rect 352 -125 353 -124
rect 353 -125 354 -124
rect 354 -125 355 -124
rect 355 -125 356 -124
rect 356 -125 357 -124
rect 357 -125 358 -124
rect 358 -125 359 -124
rect 359 -125 360 -124
rect 360 -125 361 -124
rect 361 -125 362 -124
rect 362 -125 363 -124
rect 363 -125 364 -124
rect 364 -125 365 -124
rect 365 -125 366 -124
rect 366 -125 367 -124
rect 367 -125 368 -124
rect 368 -125 369 -124
rect 369 -125 370 -124
rect 370 -125 371 -124
rect 371 -125 372 -124
rect 372 -125 373 -124
rect 373 -125 374 -124
rect 374 -125 375 -124
rect 375 -125 376 -124
rect 376 -125 377 -124
rect 377 -125 378 -124
rect 378 -125 379 -124
rect 379 -125 380 -124
rect 380 -125 381 -124
rect 381 -125 382 -124
rect 382 -125 383 -124
rect 383 -125 384 -124
rect 384 -125 385 -124
rect 385 -125 386 -124
rect 386 -125 387 -124
rect 387 -125 388 -124
rect 388 -125 389 -124
rect 389 -125 390 -124
rect 390 -125 391 -124
rect 391 -125 392 -124
rect 392 -125 393 -124
rect 393 -125 394 -124
rect 394 -125 395 -124
rect 395 -125 396 -124
rect 396 -125 397 -124
rect 397 -125 398 -124
rect 398 -125 399 -124
rect 399 -125 400 -124
rect 400 -125 401 -124
rect 401 -125 402 -124
rect 402 -125 403 -124
rect 403 -125 404 -124
rect 404 -125 405 -124
rect 405 -125 406 -124
rect 406 -125 407 -124
rect 407 -125 408 -124
rect 408 -125 409 -124
rect 409 -125 410 -124
rect 410 -125 411 -124
rect 411 -125 412 -124
rect 412 -125 413 -124
rect 413 -125 414 -124
rect 414 -125 415 -124
rect 415 -125 416 -124
rect 416 -125 417 -124
rect 417 -125 418 -124
rect 418 -125 419 -124
rect 419 -125 420 -124
rect 420 -125 421 -124
rect 421 -125 422 -124
rect 422 -125 423 -124
rect 423 -125 424 -124
rect 424 -125 425 -124
rect 425 -125 426 -124
rect 426 -125 427 -124
rect 427 -125 428 -124
rect 428 -125 429 -124
rect 429 -125 430 -124
rect 430 -125 431 -124
rect 431 -125 432 -124
rect 432 -125 433 -124
rect 433 -125 434 -124
rect 434 -125 435 -124
rect 435 -125 436 -124
rect 436 -125 437 -124
rect 437 -125 438 -124
rect 438 -125 439 -124
rect 439 -125 440 -124
rect 440 -125 441 -124
rect 441 -125 442 -124
rect 442 -125 443 -124
rect 443 -125 444 -124
rect 444 -125 445 -124
rect 445 -125 446 -124
rect 446 -125 447 -124
rect 447 -125 448 -124
rect 448 -125 449 -124
rect 449 -125 450 -124
rect 450 -125 451 -124
rect 451 -125 452 -124
rect 452 -125 453 -124
rect 453 -125 454 -124
rect 454 -125 455 -124
rect 455 -125 456 -124
rect 456 -125 457 -124
rect 457 -125 458 -124
rect 458 -125 459 -124
rect 459 -125 460 -124
rect 460 -125 461 -124
rect 461 -125 462 -124
rect 462 -125 463 -124
rect 463 -125 464 -124
rect 464 -125 465 -124
rect 465 -125 466 -124
rect 466 -125 467 -124
rect 467 -125 468 -124
rect 468 -125 469 -124
rect 469 -125 470 -124
rect 470 -125 471 -124
rect 471 -125 472 -124
rect 472 -125 473 -124
rect 473 -125 474 -124
rect 474 -125 475 -124
rect 475 -125 476 -124
rect 476 -125 477 -124
rect 477 -125 478 -124
rect 478 -125 479 -124
rect 479 -125 480 -124
rect 2 -126 3 -125
rect 3 -126 4 -125
rect 4 -126 5 -125
rect 5 -126 6 -125
rect 6 -126 7 -125
rect 7 -126 8 -125
rect 8 -126 9 -125
rect 9 -126 10 -125
rect 10 -126 11 -125
rect 11 -126 12 -125
rect 21 -126 22 -125
rect 22 -126 23 -125
rect 23 -126 24 -125
rect 24 -126 25 -125
rect 25 -126 26 -125
rect 26 -126 27 -125
rect 27 -126 28 -125
rect 28 -126 29 -125
rect 29 -126 30 -125
rect 30 -126 31 -125
rect 31 -126 32 -125
rect 32 -126 33 -125
rect 33 -126 34 -125
rect 34 -126 35 -125
rect 35 -126 36 -125
rect 36 -126 37 -125
rect 37 -126 38 -125
rect 38 -126 39 -125
rect 39 -126 40 -125
rect 40 -126 41 -125
rect 41 -126 42 -125
rect 42 -126 43 -125
rect 43 -126 44 -125
rect 53 -126 54 -125
rect 54 -126 55 -125
rect 55 -126 56 -125
rect 56 -126 57 -125
rect 57 -126 58 -125
rect 58 -126 59 -125
rect 59 -126 60 -125
rect 60 -126 61 -125
rect 61 -126 62 -125
rect 62 -126 63 -125
rect 63 -126 64 -125
rect 64 -126 65 -125
rect 65 -126 66 -125
rect 66 -126 67 -125
rect 67 -126 68 -125
rect 68 -126 69 -125
rect 69 -126 70 -125
rect 70 -126 71 -125
rect 71 -126 72 -125
rect 72 -126 73 -125
rect 73 -126 74 -125
rect 74 -126 75 -125
rect 75 -126 76 -125
rect 85 -126 86 -125
rect 86 -126 87 -125
rect 87 -126 88 -125
rect 88 -126 89 -125
rect 89 -126 90 -125
rect 90 -126 91 -125
rect 91 -126 92 -125
rect 92 -126 93 -125
rect 93 -126 94 -125
rect 94 -126 95 -125
rect 95 -126 96 -125
rect 96 -126 97 -125
rect 97 -126 98 -125
rect 98 -126 99 -125
rect 99 -126 100 -125
rect 100 -126 101 -125
rect 101 -126 102 -125
rect 102 -126 103 -125
rect 103 -126 104 -125
rect 104 -126 105 -125
rect 105 -126 106 -125
rect 106 -126 107 -125
rect 107 -126 108 -125
rect 117 -126 118 -125
rect 118 -126 119 -125
rect 119 -126 120 -125
rect 120 -126 121 -125
rect 121 -126 122 -125
rect 122 -126 123 -125
rect 123 -126 124 -125
rect 124 -126 125 -125
rect 125 -126 126 -125
rect 126 -126 127 -125
rect 127 -126 128 -125
rect 128 -126 129 -125
rect 129 -126 130 -125
rect 130 -126 131 -125
rect 131 -126 132 -125
rect 132 -126 133 -125
rect 133 -126 134 -125
rect 134 -126 135 -125
rect 135 -126 136 -125
rect 136 -126 137 -125
rect 137 -126 138 -125
rect 138 -126 139 -125
rect 139 -126 140 -125
rect 149 -126 150 -125
rect 150 -126 151 -125
rect 151 -126 152 -125
rect 152 -126 153 -125
rect 153 -126 154 -125
rect 154 -126 155 -125
rect 155 -126 156 -125
rect 156 -126 157 -125
rect 157 -126 158 -125
rect 158 -126 159 -125
rect 159 -126 160 -125
rect 160 -126 161 -125
rect 161 -126 162 -125
rect 162 -126 163 -125
rect 163 -126 164 -125
rect 164 -126 165 -125
rect 165 -126 166 -125
rect 166 -126 167 -125
rect 167 -126 168 -125
rect 168 -126 169 -125
rect 169 -126 170 -125
rect 170 -126 171 -125
rect 171 -126 172 -125
rect 181 -126 182 -125
rect 182 -126 183 -125
rect 183 -126 184 -125
rect 184 -126 185 -125
rect 185 -126 186 -125
rect 186 -126 187 -125
rect 187 -126 188 -125
rect 188 -126 189 -125
rect 189 -126 190 -125
rect 190 -126 191 -125
rect 191 -126 192 -125
rect 192 -126 193 -125
rect 193 -126 194 -125
rect 194 -126 195 -125
rect 195 -126 196 -125
rect 196 -126 197 -125
rect 197 -126 198 -125
rect 198 -126 199 -125
rect 199 -126 200 -125
rect 200 -126 201 -125
rect 201 -126 202 -125
rect 202 -126 203 -125
rect 203 -126 204 -125
rect 204 -126 205 -125
rect 205 -126 206 -125
rect 206 -126 207 -125
rect 207 -126 208 -125
rect 208 -126 209 -125
rect 209 -126 210 -125
rect 210 -126 211 -125
rect 211 -126 212 -125
rect 212 -126 213 -125
rect 213 -126 214 -125
rect 214 -126 215 -125
rect 215 -126 216 -125
rect 216 -126 217 -125
rect 217 -126 218 -125
rect 218 -126 219 -125
rect 219 -126 220 -125
rect 220 -126 221 -125
rect 221 -126 222 -125
rect 222 -126 223 -125
rect 223 -126 224 -125
rect 224 -126 225 -125
rect 225 -126 226 -125
rect 226 -126 227 -125
rect 227 -126 228 -125
rect 228 -126 229 -125
rect 229 -126 230 -125
rect 230 -126 231 -125
rect 231 -126 232 -125
rect 232 -126 233 -125
rect 233 -126 234 -125
rect 234 -126 235 -125
rect 235 -126 236 -125
rect 236 -126 237 -125
rect 237 -126 238 -125
rect 238 -126 239 -125
rect 239 -126 240 -125
rect 240 -126 241 -125
rect 241 -126 242 -125
rect 242 -126 243 -125
rect 243 -126 244 -125
rect 244 -126 245 -125
rect 245 -126 246 -125
rect 246 -126 247 -125
rect 247 -126 248 -125
rect 248 -126 249 -125
rect 249 -126 250 -125
rect 250 -126 251 -125
rect 251 -126 252 -125
rect 252 -126 253 -125
rect 253 -126 254 -125
rect 254 -126 255 -125
rect 255 -126 256 -125
rect 256 -126 257 -125
rect 257 -126 258 -125
rect 258 -126 259 -125
rect 259 -126 260 -125
rect 260 -126 261 -125
rect 261 -126 262 -125
rect 262 -126 263 -125
rect 263 -126 264 -125
rect 264 -126 265 -125
rect 265 -126 266 -125
rect 266 -126 267 -125
rect 267 -126 268 -125
rect 268 -126 269 -125
rect 269 -126 270 -125
rect 270 -126 271 -125
rect 271 -126 272 -125
rect 272 -126 273 -125
rect 273 -126 274 -125
rect 274 -126 275 -125
rect 275 -126 276 -125
rect 276 -126 277 -125
rect 277 -126 278 -125
rect 278 -126 279 -125
rect 279 -126 280 -125
rect 280 -126 281 -125
rect 281 -126 282 -125
rect 282 -126 283 -125
rect 283 -126 284 -125
rect 284 -126 285 -125
rect 285 -126 286 -125
rect 286 -126 287 -125
rect 287 -126 288 -125
rect 288 -126 289 -125
rect 289 -126 290 -125
rect 290 -126 291 -125
rect 291 -126 292 -125
rect 292 -126 293 -125
rect 293 -126 294 -125
rect 294 -126 295 -125
rect 295 -126 296 -125
rect 296 -126 297 -125
rect 297 -126 298 -125
rect 298 -126 299 -125
rect 299 -126 300 -125
rect 300 -126 301 -125
rect 301 -126 302 -125
rect 302 -126 303 -125
rect 303 -126 304 -125
rect 304 -126 305 -125
rect 305 -126 306 -125
rect 306 -126 307 -125
rect 307 -126 308 -125
rect 308 -126 309 -125
rect 309 -126 310 -125
rect 310 -126 311 -125
rect 311 -126 312 -125
rect 312 -126 313 -125
rect 313 -126 314 -125
rect 314 -126 315 -125
rect 315 -126 316 -125
rect 316 -126 317 -125
rect 317 -126 318 -125
rect 318 -126 319 -125
rect 319 -126 320 -125
rect 320 -126 321 -125
rect 321 -126 322 -125
rect 322 -126 323 -125
rect 323 -126 324 -125
rect 324 -126 325 -125
rect 325 -126 326 -125
rect 326 -126 327 -125
rect 327 -126 328 -125
rect 328 -126 329 -125
rect 329 -126 330 -125
rect 330 -126 331 -125
rect 331 -126 332 -125
rect 332 -126 333 -125
rect 333 -126 334 -125
rect 334 -126 335 -125
rect 335 -126 336 -125
rect 336 -126 337 -125
rect 337 -126 338 -125
rect 338 -126 339 -125
rect 339 -126 340 -125
rect 340 -126 341 -125
rect 341 -126 342 -125
rect 342 -126 343 -125
rect 343 -126 344 -125
rect 344 -126 345 -125
rect 345 -126 346 -125
rect 346 -126 347 -125
rect 347 -126 348 -125
rect 348 -126 349 -125
rect 349 -126 350 -125
rect 350 -126 351 -125
rect 351 -126 352 -125
rect 352 -126 353 -125
rect 353 -126 354 -125
rect 354 -126 355 -125
rect 355 -126 356 -125
rect 356 -126 357 -125
rect 357 -126 358 -125
rect 358 -126 359 -125
rect 359 -126 360 -125
rect 360 -126 361 -125
rect 361 -126 362 -125
rect 362 -126 363 -125
rect 363 -126 364 -125
rect 364 -126 365 -125
rect 365 -126 366 -125
rect 366 -126 367 -125
rect 367 -126 368 -125
rect 368 -126 369 -125
rect 369 -126 370 -125
rect 370 -126 371 -125
rect 371 -126 372 -125
rect 372 -126 373 -125
rect 373 -126 374 -125
rect 374 -126 375 -125
rect 375 -126 376 -125
rect 376 -126 377 -125
rect 377 -126 378 -125
rect 378 -126 379 -125
rect 379 -126 380 -125
rect 380 -126 381 -125
rect 381 -126 382 -125
rect 382 -126 383 -125
rect 383 -126 384 -125
rect 384 -126 385 -125
rect 385 -126 386 -125
rect 386 -126 387 -125
rect 387 -126 388 -125
rect 388 -126 389 -125
rect 389 -126 390 -125
rect 390 -126 391 -125
rect 391 -126 392 -125
rect 392 -126 393 -125
rect 393 -126 394 -125
rect 394 -126 395 -125
rect 395 -126 396 -125
rect 396 -126 397 -125
rect 397 -126 398 -125
rect 398 -126 399 -125
rect 399 -126 400 -125
rect 400 -126 401 -125
rect 401 -126 402 -125
rect 402 -126 403 -125
rect 403 -126 404 -125
rect 404 -126 405 -125
rect 405 -126 406 -125
rect 406 -126 407 -125
rect 407 -126 408 -125
rect 408 -126 409 -125
rect 409 -126 410 -125
rect 410 -126 411 -125
rect 411 -126 412 -125
rect 412 -126 413 -125
rect 413 -126 414 -125
rect 414 -126 415 -125
rect 415 -126 416 -125
rect 416 -126 417 -125
rect 417 -126 418 -125
rect 418 -126 419 -125
rect 419 -126 420 -125
rect 420 -126 421 -125
rect 421 -126 422 -125
rect 422 -126 423 -125
rect 423 -126 424 -125
rect 424 -126 425 -125
rect 425 -126 426 -125
rect 426 -126 427 -125
rect 427 -126 428 -125
rect 428 -126 429 -125
rect 429 -126 430 -125
rect 430 -126 431 -125
rect 431 -126 432 -125
rect 432 -126 433 -125
rect 433 -126 434 -125
rect 434 -126 435 -125
rect 435 -126 436 -125
rect 436 -126 437 -125
rect 437 -126 438 -125
rect 438 -126 439 -125
rect 439 -126 440 -125
rect 440 -126 441 -125
rect 441 -126 442 -125
rect 442 -126 443 -125
rect 443 -126 444 -125
rect 444 -126 445 -125
rect 445 -126 446 -125
rect 446 -126 447 -125
rect 447 -126 448 -125
rect 448 -126 449 -125
rect 449 -126 450 -125
rect 450 -126 451 -125
rect 451 -126 452 -125
rect 452 -126 453 -125
rect 453 -126 454 -125
rect 454 -126 455 -125
rect 455 -126 456 -125
rect 456 -126 457 -125
rect 457 -126 458 -125
rect 458 -126 459 -125
rect 459 -126 460 -125
rect 460 -126 461 -125
rect 461 -126 462 -125
rect 462 -126 463 -125
rect 463 -126 464 -125
rect 464 -126 465 -125
rect 465 -126 466 -125
rect 466 -126 467 -125
rect 467 -126 468 -125
rect 468 -126 469 -125
rect 469 -126 470 -125
rect 470 -126 471 -125
rect 471 -126 472 -125
rect 472 -126 473 -125
rect 473 -126 474 -125
rect 474 -126 475 -125
rect 475 -126 476 -125
rect 476 -126 477 -125
rect 477 -126 478 -125
rect 478 -126 479 -125
rect 479 -126 480 -125
rect 2 -127 3 -126
rect 3 -127 4 -126
rect 4 -127 5 -126
rect 5 -127 6 -126
rect 6 -127 7 -126
rect 7 -127 8 -126
rect 8 -127 9 -126
rect 9 -127 10 -126
rect 10 -127 11 -126
rect 11 -127 12 -126
rect 16 -127 17 -126
rect 17 -127 18 -126
rect 22 -127 23 -126
rect 23 -127 24 -126
rect 24 -127 25 -126
rect 25 -127 26 -126
rect 26 -127 27 -126
rect 27 -127 28 -126
rect 28 -127 29 -126
rect 29 -127 30 -126
rect 30 -127 31 -126
rect 31 -127 32 -126
rect 32 -127 33 -126
rect 33 -127 34 -126
rect 34 -127 35 -126
rect 35 -127 36 -126
rect 36 -127 37 -126
rect 37 -127 38 -126
rect 38 -127 39 -126
rect 39 -127 40 -126
rect 40 -127 41 -126
rect 41 -127 42 -126
rect 42 -127 43 -126
rect 43 -127 44 -126
rect 48 -127 49 -126
rect 49 -127 50 -126
rect 54 -127 55 -126
rect 55 -127 56 -126
rect 56 -127 57 -126
rect 57 -127 58 -126
rect 58 -127 59 -126
rect 59 -127 60 -126
rect 60 -127 61 -126
rect 61 -127 62 -126
rect 62 -127 63 -126
rect 63 -127 64 -126
rect 64 -127 65 -126
rect 65 -127 66 -126
rect 66 -127 67 -126
rect 67 -127 68 -126
rect 68 -127 69 -126
rect 69 -127 70 -126
rect 70 -127 71 -126
rect 71 -127 72 -126
rect 72 -127 73 -126
rect 73 -127 74 -126
rect 74 -127 75 -126
rect 75 -127 76 -126
rect 80 -127 81 -126
rect 81 -127 82 -126
rect 86 -127 87 -126
rect 87 -127 88 -126
rect 88 -127 89 -126
rect 89 -127 90 -126
rect 90 -127 91 -126
rect 91 -127 92 -126
rect 92 -127 93 -126
rect 93 -127 94 -126
rect 94 -127 95 -126
rect 95 -127 96 -126
rect 96 -127 97 -126
rect 97 -127 98 -126
rect 98 -127 99 -126
rect 99 -127 100 -126
rect 100 -127 101 -126
rect 101 -127 102 -126
rect 102 -127 103 -126
rect 103 -127 104 -126
rect 104 -127 105 -126
rect 105 -127 106 -126
rect 106 -127 107 -126
rect 107 -127 108 -126
rect 112 -127 113 -126
rect 113 -127 114 -126
rect 118 -127 119 -126
rect 119 -127 120 -126
rect 120 -127 121 -126
rect 121 -127 122 -126
rect 122 -127 123 -126
rect 123 -127 124 -126
rect 124 -127 125 -126
rect 125 -127 126 -126
rect 126 -127 127 -126
rect 127 -127 128 -126
rect 128 -127 129 -126
rect 129 -127 130 -126
rect 130 -127 131 -126
rect 131 -127 132 -126
rect 132 -127 133 -126
rect 133 -127 134 -126
rect 134 -127 135 -126
rect 135 -127 136 -126
rect 136 -127 137 -126
rect 137 -127 138 -126
rect 138 -127 139 -126
rect 139 -127 140 -126
rect 144 -127 145 -126
rect 145 -127 146 -126
rect 150 -127 151 -126
rect 151 -127 152 -126
rect 152 -127 153 -126
rect 153 -127 154 -126
rect 154 -127 155 -126
rect 155 -127 156 -126
rect 156 -127 157 -126
rect 157 -127 158 -126
rect 158 -127 159 -126
rect 159 -127 160 -126
rect 160 -127 161 -126
rect 161 -127 162 -126
rect 162 -127 163 -126
rect 163 -127 164 -126
rect 164 -127 165 -126
rect 165 -127 166 -126
rect 166 -127 167 -126
rect 167 -127 168 -126
rect 168 -127 169 -126
rect 169 -127 170 -126
rect 170 -127 171 -126
rect 171 -127 172 -126
rect 176 -127 177 -126
rect 177 -127 178 -126
rect 182 -127 183 -126
rect 183 -127 184 -126
rect 184 -127 185 -126
rect 185 -127 186 -126
rect 186 -127 187 -126
rect 187 -127 188 -126
rect 188 -127 189 -126
rect 189 -127 190 -126
rect 190 -127 191 -126
rect 191 -127 192 -126
rect 192 -127 193 -126
rect 193 -127 194 -126
rect 194 -127 195 -126
rect 195 -127 196 -126
rect 196 -127 197 -126
rect 197 -127 198 -126
rect 198 -127 199 -126
rect 199 -127 200 -126
rect 200 -127 201 -126
rect 201 -127 202 -126
rect 202 -127 203 -126
rect 203 -127 204 -126
rect 204 -127 205 -126
rect 205 -127 206 -126
rect 206 -127 207 -126
rect 207 -127 208 -126
rect 208 -127 209 -126
rect 209 -127 210 -126
rect 210 -127 211 -126
rect 211 -127 212 -126
rect 212 -127 213 -126
rect 213 -127 214 -126
rect 214 -127 215 -126
rect 215 -127 216 -126
rect 216 -127 217 -126
rect 217 -127 218 -126
rect 218 -127 219 -126
rect 219 -127 220 -126
rect 220 -127 221 -126
rect 221 -127 222 -126
rect 222 -127 223 -126
rect 223 -127 224 -126
rect 224 -127 225 -126
rect 225 -127 226 -126
rect 226 -127 227 -126
rect 227 -127 228 -126
rect 228 -127 229 -126
rect 229 -127 230 -126
rect 230 -127 231 -126
rect 231 -127 232 -126
rect 232 -127 233 -126
rect 233 -127 234 -126
rect 234 -127 235 -126
rect 235 -127 236 -126
rect 236 -127 237 -126
rect 237 -127 238 -126
rect 238 -127 239 -126
rect 239 -127 240 -126
rect 240 -127 241 -126
rect 241 -127 242 -126
rect 242 -127 243 -126
rect 243 -127 244 -126
rect 244 -127 245 -126
rect 245 -127 246 -126
rect 246 -127 247 -126
rect 247 -127 248 -126
rect 248 -127 249 -126
rect 249 -127 250 -126
rect 250 -127 251 -126
rect 251 -127 252 -126
rect 252 -127 253 -126
rect 253 -127 254 -126
rect 254 -127 255 -126
rect 255 -127 256 -126
rect 256 -127 257 -126
rect 257 -127 258 -126
rect 258 -127 259 -126
rect 259 -127 260 -126
rect 260 -127 261 -126
rect 261 -127 262 -126
rect 262 -127 263 -126
rect 263 -127 264 -126
rect 264 -127 265 -126
rect 265 -127 266 -126
rect 266 -127 267 -126
rect 267 -127 268 -126
rect 268 -127 269 -126
rect 269 -127 270 -126
rect 270 -127 271 -126
rect 271 -127 272 -126
rect 272 -127 273 -126
rect 273 -127 274 -126
rect 274 -127 275 -126
rect 275 -127 276 -126
rect 276 -127 277 -126
rect 277 -127 278 -126
rect 278 -127 279 -126
rect 279 -127 280 -126
rect 280 -127 281 -126
rect 281 -127 282 -126
rect 282 -127 283 -126
rect 283 -127 284 -126
rect 284 -127 285 -126
rect 285 -127 286 -126
rect 286 -127 287 -126
rect 287 -127 288 -126
rect 288 -127 289 -126
rect 289 -127 290 -126
rect 290 -127 291 -126
rect 291 -127 292 -126
rect 292 -127 293 -126
rect 293 -127 294 -126
rect 294 -127 295 -126
rect 295 -127 296 -126
rect 296 -127 297 -126
rect 297 -127 298 -126
rect 298 -127 299 -126
rect 299 -127 300 -126
rect 300 -127 301 -126
rect 301 -127 302 -126
rect 302 -127 303 -126
rect 303 -127 304 -126
rect 304 -127 305 -126
rect 305 -127 306 -126
rect 306 -127 307 -126
rect 307 -127 308 -126
rect 308 -127 309 -126
rect 309 -127 310 -126
rect 310 -127 311 -126
rect 311 -127 312 -126
rect 312 -127 313 -126
rect 313 -127 314 -126
rect 314 -127 315 -126
rect 315 -127 316 -126
rect 316 -127 317 -126
rect 317 -127 318 -126
rect 318 -127 319 -126
rect 319 -127 320 -126
rect 320 -127 321 -126
rect 321 -127 322 -126
rect 322 -127 323 -126
rect 323 -127 324 -126
rect 324 -127 325 -126
rect 325 -127 326 -126
rect 326 -127 327 -126
rect 327 -127 328 -126
rect 328 -127 329 -126
rect 329 -127 330 -126
rect 330 -127 331 -126
rect 331 -127 332 -126
rect 332 -127 333 -126
rect 333 -127 334 -126
rect 334 -127 335 -126
rect 335 -127 336 -126
rect 336 -127 337 -126
rect 337 -127 338 -126
rect 338 -127 339 -126
rect 339 -127 340 -126
rect 340 -127 341 -126
rect 341 -127 342 -126
rect 342 -127 343 -126
rect 343 -127 344 -126
rect 344 -127 345 -126
rect 345 -127 346 -126
rect 346 -127 347 -126
rect 347 -127 348 -126
rect 348 -127 349 -126
rect 349 -127 350 -126
rect 350 -127 351 -126
rect 351 -127 352 -126
rect 352 -127 353 -126
rect 353 -127 354 -126
rect 354 -127 355 -126
rect 355 -127 356 -126
rect 356 -127 357 -126
rect 357 -127 358 -126
rect 358 -127 359 -126
rect 359 -127 360 -126
rect 360 -127 361 -126
rect 361 -127 362 -126
rect 362 -127 363 -126
rect 363 -127 364 -126
rect 364 -127 365 -126
rect 365 -127 366 -126
rect 366 -127 367 -126
rect 367 -127 368 -126
rect 368 -127 369 -126
rect 369 -127 370 -126
rect 370 -127 371 -126
rect 371 -127 372 -126
rect 372 -127 373 -126
rect 373 -127 374 -126
rect 374 -127 375 -126
rect 375 -127 376 -126
rect 376 -127 377 -126
rect 377 -127 378 -126
rect 378 -127 379 -126
rect 379 -127 380 -126
rect 380 -127 381 -126
rect 381 -127 382 -126
rect 382 -127 383 -126
rect 383 -127 384 -126
rect 384 -127 385 -126
rect 385 -127 386 -126
rect 386 -127 387 -126
rect 387 -127 388 -126
rect 388 -127 389 -126
rect 389 -127 390 -126
rect 390 -127 391 -126
rect 391 -127 392 -126
rect 392 -127 393 -126
rect 393 -127 394 -126
rect 394 -127 395 -126
rect 395 -127 396 -126
rect 396 -127 397 -126
rect 397 -127 398 -126
rect 398 -127 399 -126
rect 399 -127 400 -126
rect 400 -127 401 -126
rect 401 -127 402 -126
rect 402 -127 403 -126
rect 403 -127 404 -126
rect 404 -127 405 -126
rect 405 -127 406 -126
rect 406 -127 407 -126
rect 407 -127 408 -126
rect 408 -127 409 -126
rect 409 -127 410 -126
rect 410 -127 411 -126
rect 411 -127 412 -126
rect 412 -127 413 -126
rect 413 -127 414 -126
rect 414 -127 415 -126
rect 415 -127 416 -126
rect 416 -127 417 -126
rect 417 -127 418 -126
rect 418 -127 419 -126
rect 419 -127 420 -126
rect 420 -127 421 -126
rect 421 -127 422 -126
rect 422 -127 423 -126
rect 423 -127 424 -126
rect 424 -127 425 -126
rect 425 -127 426 -126
rect 426 -127 427 -126
rect 427 -127 428 -126
rect 428 -127 429 -126
rect 429 -127 430 -126
rect 430 -127 431 -126
rect 431 -127 432 -126
rect 432 -127 433 -126
rect 433 -127 434 -126
rect 434 -127 435 -126
rect 435 -127 436 -126
rect 436 -127 437 -126
rect 437 -127 438 -126
rect 438 -127 439 -126
rect 439 -127 440 -126
rect 440 -127 441 -126
rect 441 -127 442 -126
rect 442 -127 443 -126
rect 443 -127 444 -126
rect 444 -127 445 -126
rect 445 -127 446 -126
rect 446 -127 447 -126
rect 447 -127 448 -126
rect 448 -127 449 -126
rect 449 -127 450 -126
rect 450 -127 451 -126
rect 451 -127 452 -126
rect 452 -127 453 -126
rect 453 -127 454 -126
rect 454 -127 455 -126
rect 455 -127 456 -126
rect 456 -127 457 -126
rect 457 -127 458 -126
rect 458 -127 459 -126
rect 459 -127 460 -126
rect 460 -127 461 -126
rect 461 -127 462 -126
rect 462 -127 463 -126
rect 463 -127 464 -126
rect 464 -127 465 -126
rect 465 -127 466 -126
rect 466 -127 467 -126
rect 467 -127 468 -126
rect 468 -127 469 -126
rect 469 -127 470 -126
rect 470 -127 471 -126
rect 471 -127 472 -126
rect 472 -127 473 -126
rect 473 -127 474 -126
rect 474 -127 475 -126
rect 475 -127 476 -126
rect 476 -127 477 -126
rect 477 -127 478 -126
rect 478 -127 479 -126
rect 479 -127 480 -126
rect 2 -128 3 -127
rect 3 -128 4 -127
rect 4 -128 5 -127
rect 5 -128 6 -127
rect 6 -128 7 -127
rect 7 -128 8 -127
rect 8 -128 9 -127
rect 9 -128 10 -127
rect 10 -128 11 -127
rect 11 -128 12 -127
rect 15 -128 16 -127
rect 16 -128 17 -127
rect 17 -128 18 -127
rect 18 -128 19 -127
rect 22 -128 23 -127
rect 23 -128 24 -127
rect 24 -128 25 -127
rect 25 -128 26 -127
rect 26 -128 27 -127
rect 27 -128 28 -127
rect 28 -128 29 -127
rect 29 -128 30 -127
rect 30 -128 31 -127
rect 31 -128 32 -127
rect 32 -128 33 -127
rect 33 -128 34 -127
rect 34 -128 35 -127
rect 35 -128 36 -127
rect 36 -128 37 -127
rect 37 -128 38 -127
rect 38 -128 39 -127
rect 39 -128 40 -127
rect 40 -128 41 -127
rect 41 -128 42 -127
rect 42 -128 43 -127
rect 43 -128 44 -127
rect 47 -128 48 -127
rect 48 -128 49 -127
rect 49 -128 50 -127
rect 50 -128 51 -127
rect 54 -128 55 -127
rect 55 -128 56 -127
rect 56 -128 57 -127
rect 57 -128 58 -127
rect 58 -128 59 -127
rect 59 -128 60 -127
rect 60 -128 61 -127
rect 61 -128 62 -127
rect 62 -128 63 -127
rect 63 -128 64 -127
rect 64 -128 65 -127
rect 65 -128 66 -127
rect 66 -128 67 -127
rect 67 -128 68 -127
rect 68 -128 69 -127
rect 69 -128 70 -127
rect 70 -128 71 -127
rect 71 -128 72 -127
rect 72 -128 73 -127
rect 73 -128 74 -127
rect 74 -128 75 -127
rect 75 -128 76 -127
rect 79 -128 80 -127
rect 80 -128 81 -127
rect 81 -128 82 -127
rect 82 -128 83 -127
rect 86 -128 87 -127
rect 87 -128 88 -127
rect 88 -128 89 -127
rect 89 -128 90 -127
rect 90 -128 91 -127
rect 91 -128 92 -127
rect 92 -128 93 -127
rect 93 -128 94 -127
rect 94 -128 95 -127
rect 95 -128 96 -127
rect 96 -128 97 -127
rect 97 -128 98 -127
rect 98 -128 99 -127
rect 99 -128 100 -127
rect 100 -128 101 -127
rect 101 -128 102 -127
rect 102 -128 103 -127
rect 103 -128 104 -127
rect 104 -128 105 -127
rect 105 -128 106 -127
rect 106 -128 107 -127
rect 107 -128 108 -127
rect 111 -128 112 -127
rect 112 -128 113 -127
rect 113 -128 114 -127
rect 114 -128 115 -127
rect 118 -128 119 -127
rect 119 -128 120 -127
rect 120 -128 121 -127
rect 121 -128 122 -127
rect 122 -128 123 -127
rect 123 -128 124 -127
rect 124 -128 125 -127
rect 125 -128 126 -127
rect 126 -128 127 -127
rect 127 -128 128 -127
rect 128 -128 129 -127
rect 129 -128 130 -127
rect 130 -128 131 -127
rect 131 -128 132 -127
rect 132 -128 133 -127
rect 133 -128 134 -127
rect 134 -128 135 -127
rect 135 -128 136 -127
rect 136 -128 137 -127
rect 137 -128 138 -127
rect 138 -128 139 -127
rect 139 -128 140 -127
rect 143 -128 144 -127
rect 144 -128 145 -127
rect 145 -128 146 -127
rect 146 -128 147 -127
rect 150 -128 151 -127
rect 151 -128 152 -127
rect 152 -128 153 -127
rect 153 -128 154 -127
rect 154 -128 155 -127
rect 155 -128 156 -127
rect 156 -128 157 -127
rect 157 -128 158 -127
rect 158 -128 159 -127
rect 159 -128 160 -127
rect 160 -128 161 -127
rect 161 -128 162 -127
rect 162 -128 163 -127
rect 163 -128 164 -127
rect 164 -128 165 -127
rect 165 -128 166 -127
rect 166 -128 167 -127
rect 167 -128 168 -127
rect 168 -128 169 -127
rect 169 -128 170 -127
rect 170 -128 171 -127
rect 171 -128 172 -127
rect 175 -128 176 -127
rect 176 -128 177 -127
rect 177 -128 178 -127
rect 178 -128 179 -127
rect 182 -128 183 -127
rect 183 -128 184 -127
rect 184 -128 185 -127
rect 185 -128 186 -127
rect 186 -128 187 -127
rect 187 -128 188 -127
rect 188 -128 189 -127
rect 189 -128 190 -127
rect 190 -128 191 -127
rect 191 -128 192 -127
rect 192 -128 193 -127
rect 193 -128 194 -127
rect 194 -128 195 -127
rect 195 -128 196 -127
rect 196 -128 197 -127
rect 197 -128 198 -127
rect 198 -128 199 -127
rect 199 -128 200 -127
rect 200 -128 201 -127
rect 201 -128 202 -127
rect 202 -128 203 -127
rect 203 -128 204 -127
rect 204 -128 205 -127
rect 205 -128 206 -127
rect 206 -128 207 -127
rect 207 -128 208 -127
rect 208 -128 209 -127
rect 209 -128 210 -127
rect 210 -128 211 -127
rect 211 -128 212 -127
rect 212 -128 213 -127
rect 213 -128 214 -127
rect 214 -128 215 -127
rect 215 -128 216 -127
rect 216 -128 217 -127
rect 217 -128 218 -127
rect 218 -128 219 -127
rect 219 -128 220 -127
rect 220 -128 221 -127
rect 221 -128 222 -127
rect 222 -128 223 -127
rect 223 -128 224 -127
rect 224 -128 225 -127
rect 225 -128 226 -127
rect 226 -128 227 -127
rect 227 -128 228 -127
rect 228 -128 229 -127
rect 229 -128 230 -127
rect 230 -128 231 -127
rect 231 -128 232 -127
rect 232 -128 233 -127
rect 233 -128 234 -127
rect 234 -128 235 -127
rect 235 -128 236 -127
rect 236 -128 237 -127
rect 237 -128 238 -127
rect 238 -128 239 -127
rect 239 -128 240 -127
rect 240 -128 241 -127
rect 241 -128 242 -127
rect 242 -128 243 -127
rect 243 -128 244 -127
rect 244 -128 245 -127
rect 245 -128 246 -127
rect 246 -128 247 -127
rect 247 -128 248 -127
rect 248 -128 249 -127
rect 249 -128 250 -127
rect 250 -128 251 -127
rect 251 -128 252 -127
rect 252 -128 253 -127
rect 253 -128 254 -127
rect 254 -128 255 -127
rect 255 -128 256 -127
rect 256 -128 257 -127
rect 257 -128 258 -127
rect 258 -128 259 -127
rect 259 -128 260 -127
rect 260 -128 261 -127
rect 261 -128 262 -127
rect 262 -128 263 -127
rect 263 -128 264 -127
rect 264 -128 265 -127
rect 265 -128 266 -127
rect 266 -128 267 -127
rect 267 -128 268 -127
rect 268 -128 269 -127
rect 269 -128 270 -127
rect 270 -128 271 -127
rect 271 -128 272 -127
rect 272 -128 273 -127
rect 273 -128 274 -127
rect 274 -128 275 -127
rect 275 -128 276 -127
rect 276 -128 277 -127
rect 277 -128 278 -127
rect 278 -128 279 -127
rect 279 -128 280 -127
rect 280 -128 281 -127
rect 281 -128 282 -127
rect 282 -128 283 -127
rect 283 -128 284 -127
rect 284 -128 285 -127
rect 285 -128 286 -127
rect 286 -128 287 -127
rect 287 -128 288 -127
rect 288 -128 289 -127
rect 289 -128 290 -127
rect 290 -128 291 -127
rect 291 -128 292 -127
rect 292 -128 293 -127
rect 293 -128 294 -127
rect 294 -128 295 -127
rect 295 -128 296 -127
rect 296 -128 297 -127
rect 297 -128 298 -127
rect 298 -128 299 -127
rect 299 -128 300 -127
rect 300 -128 301 -127
rect 301 -128 302 -127
rect 302 -128 303 -127
rect 303 -128 304 -127
rect 304 -128 305 -127
rect 305 -128 306 -127
rect 306 -128 307 -127
rect 307 -128 308 -127
rect 308 -128 309 -127
rect 309 -128 310 -127
rect 310 -128 311 -127
rect 311 -128 312 -127
rect 312 -128 313 -127
rect 313 -128 314 -127
rect 314 -128 315 -127
rect 315 -128 316 -127
rect 316 -128 317 -127
rect 317 -128 318 -127
rect 318 -128 319 -127
rect 319 -128 320 -127
rect 320 -128 321 -127
rect 321 -128 322 -127
rect 322 -128 323 -127
rect 323 -128 324 -127
rect 324 -128 325 -127
rect 325 -128 326 -127
rect 326 -128 327 -127
rect 327 -128 328 -127
rect 328 -128 329 -127
rect 329 -128 330 -127
rect 330 -128 331 -127
rect 331 -128 332 -127
rect 332 -128 333 -127
rect 333 -128 334 -127
rect 334 -128 335 -127
rect 335 -128 336 -127
rect 336 -128 337 -127
rect 337 -128 338 -127
rect 338 -128 339 -127
rect 339 -128 340 -127
rect 340 -128 341 -127
rect 341 -128 342 -127
rect 342 -128 343 -127
rect 343 -128 344 -127
rect 344 -128 345 -127
rect 345 -128 346 -127
rect 346 -128 347 -127
rect 347 -128 348 -127
rect 348 -128 349 -127
rect 349 -128 350 -127
rect 350 -128 351 -127
rect 351 -128 352 -127
rect 352 -128 353 -127
rect 353 -128 354 -127
rect 354 -128 355 -127
rect 355 -128 356 -127
rect 356 -128 357 -127
rect 357 -128 358 -127
rect 358 -128 359 -127
rect 359 -128 360 -127
rect 360 -128 361 -127
rect 361 -128 362 -127
rect 362 -128 363 -127
rect 363 -128 364 -127
rect 364 -128 365 -127
rect 365 -128 366 -127
rect 366 -128 367 -127
rect 367 -128 368 -127
rect 368 -128 369 -127
rect 369 -128 370 -127
rect 370 -128 371 -127
rect 371 -128 372 -127
rect 372 -128 373 -127
rect 373 -128 374 -127
rect 374 -128 375 -127
rect 375 -128 376 -127
rect 376 -128 377 -127
rect 377 -128 378 -127
rect 378 -128 379 -127
rect 379 -128 380 -127
rect 380 -128 381 -127
rect 381 -128 382 -127
rect 382 -128 383 -127
rect 383 -128 384 -127
rect 384 -128 385 -127
rect 385 -128 386 -127
rect 386 -128 387 -127
rect 387 -128 388 -127
rect 388 -128 389 -127
rect 389 -128 390 -127
rect 390 -128 391 -127
rect 391 -128 392 -127
rect 392 -128 393 -127
rect 393 -128 394 -127
rect 394 -128 395 -127
rect 395 -128 396 -127
rect 396 -128 397 -127
rect 397 -128 398 -127
rect 398 -128 399 -127
rect 399 -128 400 -127
rect 400 -128 401 -127
rect 401 -128 402 -127
rect 402 -128 403 -127
rect 403 -128 404 -127
rect 404 -128 405 -127
rect 405 -128 406 -127
rect 406 -128 407 -127
rect 407 -128 408 -127
rect 408 -128 409 -127
rect 409 -128 410 -127
rect 410 -128 411 -127
rect 411 -128 412 -127
rect 412 -128 413 -127
rect 413 -128 414 -127
rect 414 -128 415 -127
rect 415 -128 416 -127
rect 416 -128 417 -127
rect 417 -128 418 -127
rect 418 -128 419 -127
rect 419 -128 420 -127
rect 420 -128 421 -127
rect 421 -128 422 -127
rect 422 -128 423 -127
rect 423 -128 424 -127
rect 424 -128 425 -127
rect 425 -128 426 -127
rect 426 -128 427 -127
rect 427 -128 428 -127
rect 428 -128 429 -127
rect 429 -128 430 -127
rect 430 -128 431 -127
rect 431 -128 432 -127
rect 432 -128 433 -127
rect 433 -128 434 -127
rect 434 -128 435 -127
rect 435 -128 436 -127
rect 436 -128 437 -127
rect 437 -128 438 -127
rect 438 -128 439 -127
rect 439 -128 440 -127
rect 440 -128 441 -127
rect 441 -128 442 -127
rect 442 -128 443 -127
rect 443 -128 444 -127
rect 444 -128 445 -127
rect 445 -128 446 -127
rect 446 -128 447 -127
rect 447 -128 448 -127
rect 448 -128 449 -127
rect 449 -128 450 -127
rect 450 -128 451 -127
rect 451 -128 452 -127
rect 452 -128 453 -127
rect 453 -128 454 -127
rect 454 -128 455 -127
rect 455 -128 456 -127
rect 456 -128 457 -127
rect 457 -128 458 -127
rect 458 -128 459 -127
rect 459 -128 460 -127
rect 460 -128 461 -127
rect 461 -128 462 -127
rect 462 -128 463 -127
rect 463 -128 464 -127
rect 464 -128 465 -127
rect 465 -128 466 -127
rect 466 -128 467 -127
rect 467 -128 468 -127
rect 468 -128 469 -127
rect 469 -128 470 -127
rect 470 -128 471 -127
rect 471 -128 472 -127
rect 472 -128 473 -127
rect 473 -128 474 -127
rect 474 -128 475 -127
rect 475 -128 476 -127
rect 476 -128 477 -127
rect 477 -128 478 -127
rect 478 -128 479 -127
rect 479 -128 480 -127
rect 2 -129 3 -128
rect 3 -129 4 -128
rect 4 -129 5 -128
rect 5 -129 6 -128
rect 6 -129 7 -128
rect 7 -129 8 -128
rect 8 -129 9 -128
rect 9 -129 10 -128
rect 10 -129 11 -128
rect 11 -129 12 -128
rect 12 -129 13 -128
rect 13 -129 14 -128
rect 14 -129 15 -128
rect 15 -129 16 -128
rect 16 -129 17 -128
rect 17 -129 18 -128
rect 18 -129 19 -128
rect 19 -129 20 -128
rect 20 -129 21 -128
rect 21 -129 22 -128
rect 22 -129 23 -128
rect 23 -129 24 -128
rect 24 -129 25 -128
rect 25 -129 26 -128
rect 26 -129 27 -128
rect 27 -129 28 -128
rect 28 -129 29 -128
rect 29 -129 30 -128
rect 30 -129 31 -128
rect 31 -129 32 -128
rect 32 -129 33 -128
rect 33 -129 34 -128
rect 34 -129 35 -128
rect 35 -129 36 -128
rect 36 -129 37 -128
rect 37 -129 38 -128
rect 38 -129 39 -128
rect 39 -129 40 -128
rect 40 -129 41 -128
rect 41 -129 42 -128
rect 42 -129 43 -128
rect 43 -129 44 -128
rect 44 -129 45 -128
rect 45 -129 46 -128
rect 46 -129 47 -128
rect 47 -129 48 -128
rect 48 -129 49 -128
rect 49 -129 50 -128
rect 50 -129 51 -128
rect 51 -129 52 -128
rect 52 -129 53 -128
rect 53 -129 54 -128
rect 54 -129 55 -128
rect 55 -129 56 -128
rect 56 -129 57 -128
rect 57 -129 58 -128
rect 58 -129 59 -128
rect 59 -129 60 -128
rect 60 -129 61 -128
rect 61 -129 62 -128
rect 62 -129 63 -128
rect 63 -129 64 -128
rect 64 -129 65 -128
rect 65 -129 66 -128
rect 66 -129 67 -128
rect 67 -129 68 -128
rect 68 -129 69 -128
rect 69 -129 70 -128
rect 70 -129 71 -128
rect 71 -129 72 -128
rect 72 -129 73 -128
rect 73 -129 74 -128
rect 74 -129 75 -128
rect 75 -129 76 -128
rect 76 -129 77 -128
rect 77 -129 78 -128
rect 78 -129 79 -128
rect 79 -129 80 -128
rect 80 -129 81 -128
rect 81 -129 82 -128
rect 82 -129 83 -128
rect 83 -129 84 -128
rect 84 -129 85 -128
rect 85 -129 86 -128
rect 86 -129 87 -128
rect 87 -129 88 -128
rect 88 -129 89 -128
rect 89 -129 90 -128
rect 90 -129 91 -128
rect 91 -129 92 -128
rect 92 -129 93 -128
rect 93 -129 94 -128
rect 94 -129 95 -128
rect 95 -129 96 -128
rect 96 -129 97 -128
rect 97 -129 98 -128
rect 98 -129 99 -128
rect 99 -129 100 -128
rect 100 -129 101 -128
rect 101 -129 102 -128
rect 102 -129 103 -128
rect 103 -129 104 -128
rect 104 -129 105 -128
rect 105 -129 106 -128
rect 106 -129 107 -128
rect 107 -129 108 -128
rect 108 -129 109 -128
rect 109 -129 110 -128
rect 110 -129 111 -128
rect 111 -129 112 -128
rect 112 -129 113 -128
rect 113 -129 114 -128
rect 114 -129 115 -128
rect 115 -129 116 -128
rect 116 -129 117 -128
rect 117 -129 118 -128
rect 118 -129 119 -128
rect 119 -129 120 -128
rect 120 -129 121 -128
rect 121 -129 122 -128
rect 122 -129 123 -128
rect 123 -129 124 -128
rect 124 -129 125 -128
rect 125 -129 126 -128
rect 126 -129 127 -128
rect 127 -129 128 -128
rect 128 -129 129 -128
rect 129 -129 130 -128
rect 130 -129 131 -128
rect 131 -129 132 -128
rect 132 -129 133 -128
rect 133 -129 134 -128
rect 134 -129 135 -128
rect 135 -129 136 -128
rect 136 -129 137 -128
rect 137 -129 138 -128
rect 138 -129 139 -128
rect 139 -129 140 -128
rect 140 -129 141 -128
rect 141 -129 142 -128
rect 142 -129 143 -128
rect 143 -129 144 -128
rect 144 -129 145 -128
rect 145 -129 146 -128
rect 146 -129 147 -128
rect 147 -129 148 -128
rect 148 -129 149 -128
rect 149 -129 150 -128
rect 150 -129 151 -128
rect 151 -129 152 -128
rect 152 -129 153 -128
rect 153 -129 154 -128
rect 154 -129 155 -128
rect 155 -129 156 -128
rect 156 -129 157 -128
rect 157 -129 158 -128
rect 158 -129 159 -128
rect 159 -129 160 -128
rect 160 -129 161 -128
rect 161 -129 162 -128
rect 162 -129 163 -128
rect 163 -129 164 -128
rect 164 -129 165 -128
rect 165 -129 166 -128
rect 166 -129 167 -128
rect 167 -129 168 -128
rect 168 -129 169 -128
rect 169 -129 170 -128
rect 170 -129 171 -128
rect 171 -129 172 -128
rect 172 -129 173 -128
rect 173 -129 174 -128
rect 174 -129 175 -128
rect 175 -129 176 -128
rect 176 -129 177 -128
rect 177 -129 178 -128
rect 178 -129 179 -128
rect 179 -129 180 -128
rect 180 -129 181 -128
rect 181 -129 182 -128
rect 182 -129 183 -128
rect 183 -129 184 -128
rect 184 -129 185 -128
rect 185 -129 186 -128
rect 186 -129 187 -128
rect 187 -129 188 -128
rect 188 -129 189 -128
rect 189 -129 190 -128
rect 190 -129 191 -128
rect 191 -129 192 -128
rect 192 -129 193 -128
rect 193 -129 194 -128
rect 194 -129 195 -128
rect 195 -129 196 -128
rect 196 -129 197 -128
rect 197 -129 198 -128
rect 198 -129 199 -128
rect 199 -129 200 -128
rect 200 -129 201 -128
rect 201 -129 202 -128
rect 202 -129 203 -128
rect 203 -129 204 -128
rect 204 -129 205 -128
rect 205 -129 206 -128
rect 206 -129 207 -128
rect 207 -129 208 -128
rect 208 -129 209 -128
rect 209 -129 210 -128
rect 210 -129 211 -128
rect 211 -129 212 -128
rect 212 -129 213 -128
rect 213 -129 214 -128
rect 214 -129 215 -128
rect 215 -129 216 -128
rect 216 -129 217 -128
rect 217 -129 218 -128
rect 218 -129 219 -128
rect 219 -129 220 -128
rect 220 -129 221 -128
rect 221 -129 222 -128
rect 222 -129 223 -128
rect 223 -129 224 -128
rect 224 -129 225 -128
rect 225 -129 226 -128
rect 226 -129 227 -128
rect 227 -129 228 -128
rect 228 -129 229 -128
rect 229 -129 230 -128
rect 230 -129 231 -128
rect 231 -129 232 -128
rect 232 -129 233 -128
rect 233 -129 234 -128
rect 234 -129 235 -128
rect 235 -129 236 -128
rect 236 -129 237 -128
rect 237 -129 238 -128
rect 238 -129 239 -128
rect 239 -129 240 -128
rect 240 -129 241 -128
rect 241 -129 242 -128
rect 242 -129 243 -128
rect 243 -129 244 -128
rect 244 -129 245 -128
rect 245 -129 246 -128
rect 246 -129 247 -128
rect 247 -129 248 -128
rect 248 -129 249 -128
rect 249 -129 250 -128
rect 250 -129 251 -128
rect 251 -129 252 -128
rect 252 -129 253 -128
rect 253 -129 254 -128
rect 254 -129 255 -128
rect 255 -129 256 -128
rect 256 -129 257 -128
rect 257 -129 258 -128
rect 258 -129 259 -128
rect 259 -129 260 -128
rect 260 -129 261 -128
rect 261 -129 262 -128
rect 262 -129 263 -128
rect 263 -129 264 -128
rect 264 -129 265 -128
rect 265 -129 266 -128
rect 266 -129 267 -128
rect 267 -129 268 -128
rect 268 -129 269 -128
rect 269 -129 270 -128
rect 270 -129 271 -128
rect 271 -129 272 -128
rect 272 -129 273 -128
rect 273 -129 274 -128
rect 274 -129 275 -128
rect 275 -129 276 -128
rect 276 -129 277 -128
rect 277 -129 278 -128
rect 278 -129 279 -128
rect 279 -129 280 -128
rect 280 -129 281 -128
rect 281 -129 282 -128
rect 282 -129 283 -128
rect 283 -129 284 -128
rect 284 -129 285 -128
rect 285 -129 286 -128
rect 286 -129 287 -128
rect 287 -129 288 -128
rect 288 -129 289 -128
rect 289 -129 290 -128
rect 290 -129 291 -128
rect 291 -129 292 -128
rect 292 -129 293 -128
rect 293 -129 294 -128
rect 294 -129 295 -128
rect 295 -129 296 -128
rect 296 -129 297 -128
rect 297 -129 298 -128
rect 298 -129 299 -128
rect 299 -129 300 -128
rect 300 -129 301 -128
rect 301 -129 302 -128
rect 302 -129 303 -128
rect 303 -129 304 -128
rect 304 -129 305 -128
rect 305 -129 306 -128
rect 306 -129 307 -128
rect 307 -129 308 -128
rect 308 -129 309 -128
rect 309 -129 310 -128
rect 310 -129 311 -128
rect 311 -129 312 -128
rect 312 -129 313 -128
rect 313 -129 314 -128
rect 314 -129 315 -128
rect 315 -129 316 -128
rect 316 -129 317 -128
rect 317 -129 318 -128
rect 318 -129 319 -128
rect 319 -129 320 -128
rect 320 -129 321 -128
rect 321 -129 322 -128
rect 322 -129 323 -128
rect 323 -129 324 -128
rect 324 -129 325 -128
rect 325 -129 326 -128
rect 326 -129 327 -128
rect 327 -129 328 -128
rect 328 -129 329 -128
rect 329 -129 330 -128
rect 330 -129 331 -128
rect 331 -129 332 -128
rect 332 -129 333 -128
rect 333 -129 334 -128
rect 334 -129 335 -128
rect 335 -129 336 -128
rect 336 -129 337 -128
rect 337 -129 338 -128
rect 338 -129 339 -128
rect 339 -129 340 -128
rect 340 -129 341 -128
rect 341 -129 342 -128
rect 342 -129 343 -128
rect 343 -129 344 -128
rect 344 -129 345 -128
rect 345 -129 346 -128
rect 346 -129 347 -128
rect 347 -129 348 -128
rect 348 -129 349 -128
rect 349 -129 350 -128
rect 350 -129 351 -128
rect 351 -129 352 -128
rect 352 -129 353 -128
rect 353 -129 354 -128
rect 354 -129 355 -128
rect 355 -129 356 -128
rect 356 -129 357 -128
rect 357 -129 358 -128
rect 358 -129 359 -128
rect 359 -129 360 -128
rect 360 -129 361 -128
rect 361 -129 362 -128
rect 362 -129 363 -128
rect 363 -129 364 -128
rect 364 -129 365 -128
rect 365 -129 366 -128
rect 366 -129 367 -128
rect 367 -129 368 -128
rect 368 -129 369 -128
rect 369 -129 370 -128
rect 370 -129 371 -128
rect 371 -129 372 -128
rect 372 -129 373 -128
rect 373 -129 374 -128
rect 374 -129 375 -128
rect 375 -129 376 -128
rect 376 -129 377 -128
rect 377 -129 378 -128
rect 378 -129 379 -128
rect 379 -129 380 -128
rect 380 -129 381 -128
rect 381 -129 382 -128
rect 382 -129 383 -128
rect 383 -129 384 -128
rect 384 -129 385 -128
rect 385 -129 386 -128
rect 386 -129 387 -128
rect 387 -129 388 -128
rect 388 -129 389 -128
rect 389 -129 390 -128
rect 390 -129 391 -128
rect 391 -129 392 -128
rect 392 -129 393 -128
rect 393 -129 394 -128
rect 394 -129 395 -128
rect 395 -129 396 -128
rect 396 -129 397 -128
rect 397 -129 398 -128
rect 398 -129 399 -128
rect 399 -129 400 -128
rect 400 -129 401 -128
rect 401 -129 402 -128
rect 402 -129 403 -128
rect 403 -129 404 -128
rect 404 -129 405 -128
rect 405 -129 406 -128
rect 406 -129 407 -128
rect 407 -129 408 -128
rect 408 -129 409 -128
rect 409 -129 410 -128
rect 410 -129 411 -128
rect 411 -129 412 -128
rect 412 -129 413 -128
rect 413 -129 414 -128
rect 414 -129 415 -128
rect 415 -129 416 -128
rect 416 -129 417 -128
rect 417 -129 418 -128
rect 418 -129 419 -128
rect 419 -129 420 -128
rect 420 -129 421 -128
rect 421 -129 422 -128
rect 422 -129 423 -128
rect 423 -129 424 -128
rect 424 -129 425 -128
rect 425 -129 426 -128
rect 426 -129 427 -128
rect 427 -129 428 -128
rect 428 -129 429 -128
rect 429 -129 430 -128
rect 430 -129 431 -128
rect 431 -129 432 -128
rect 432 -129 433 -128
rect 433 -129 434 -128
rect 434 -129 435 -128
rect 435 -129 436 -128
rect 436 -129 437 -128
rect 437 -129 438 -128
rect 438 -129 439 -128
rect 439 -129 440 -128
rect 440 -129 441 -128
rect 441 -129 442 -128
rect 442 -129 443 -128
rect 443 -129 444 -128
rect 444 -129 445 -128
rect 445 -129 446 -128
rect 446 -129 447 -128
rect 447 -129 448 -128
rect 448 -129 449 -128
rect 449 -129 450 -128
rect 450 -129 451 -128
rect 451 -129 452 -128
rect 452 -129 453 -128
rect 453 -129 454 -128
rect 454 -129 455 -128
rect 455 -129 456 -128
rect 456 -129 457 -128
rect 457 -129 458 -128
rect 458 -129 459 -128
rect 459 -129 460 -128
rect 460 -129 461 -128
rect 461 -129 462 -128
rect 462 -129 463 -128
rect 463 -129 464 -128
rect 464 -129 465 -128
rect 465 -129 466 -128
rect 466 -129 467 -128
rect 467 -129 468 -128
rect 468 -129 469 -128
rect 469 -129 470 -128
rect 470 -129 471 -128
rect 471 -129 472 -128
rect 472 -129 473 -128
rect 473 -129 474 -128
rect 474 -129 475 -128
rect 475 -129 476 -128
rect 476 -129 477 -128
rect 477 -129 478 -128
rect 478 -129 479 -128
rect 479 -129 480 -128
rect 2 -130 3 -129
rect 3 -130 4 -129
rect 4 -130 5 -129
rect 5 -130 6 -129
rect 6 -130 7 -129
rect 7 -130 8 -129
rect 8 -130 9 -129
rect 9 -130 10 -129
rect 10 -130 11 -129
rect 11 -130 12 -129
rect 12 -130 13 -129
rect 13 -130 14 -129
rect 14 -130 15 -129
rect 15 -130 16 -129
rect 16 -130 17 -129
rect 17 -130 18 -129
rect 18 -130 19 -129
rect 19 -130 20 -129
rect 20 -130 21 -129
rect 21 -130 22 -129
rect 22 -130 23 -129
rect 23 -130 24 -129
rect 24 -130 25 -129
rect 25 -130 26 -129
rect 26 -130 27 -129
rect 27 -130 28 -129
rect 28 -130 29 -129
rect 29 -130 30 -129
rect 30 -130 31 -129
rect 31 -130 32 -129
rect 32 -130 33 -129
rect 33 -130 34 -129
rect 34 -130 35 -129
rect 35 -130 36 -129
rect 36 -130 37 -129
rect 37 -130 38 -129
rect 38 -130 39 -129
rect 39 -130 40 -129
rect 40 -130 41 -129
rect 41 -130 42 -129
rect 42 -130 43 -129
rect 43 -130 44 -129
rect 44 -130 45 -129
rect 45 -130 46 -129
rect 46 -130 47 -129
rect 47 -130 48 -129
rect 48 -130 49 -129
rect 49 -130 50 -129
rect 50 -130 51 -129
rect 51 -130 52 -129
rect 52 -130 53 -129
rect 53 -130 54 -129
rect 54 -130 55 -129
rect 55 -130 56 -129
rect 56 -130 57 -129
rect 57 -130 58 -129
rect 58 -130 59 -129
rect 59 -130 60 -129
rect 60 -130 61 -129
rect 61 -130 62 -129
rect 62 -130 63 -129
rect 63 -130 64 -129
rect 64 -130 65 -129
rect 65 -130 66 -129
rect 66 -130 67 -129
rect 67 -130 68 -129
rect 68 -130 69 -129
rect 69 -130 70 -129
rect 70 -130 71 -129
rect 71 -130 72 -129
rect 72 -130 73 -129
rect 73 -130 74 -129
rect 74 -130 75 -129
rect 75 -130 76 -129
rect 76 -130 77 -129
rect 77 -130 78 -129
rect 78 -130 79 -129
rect 79 -130 80 -129
rect 80 -130 81 -129
rect 81 -130 82 -129
rect 82 -130 83 -129
rect 83 -130 84 -129
rect 84 -130 85 -129
rect 85 -130 86 -129
rect 86 -130 87 -129
rect 87 -130 88 -129
rect 88 -130 89 -129
rect 89 -130 90 -129
rect 90 -130 91 -129
rect 91 -130 92 -129
rect 92 -130 93 -129
rect 93 -130 94 -129
rect 94 -130 95 -129
rect 95 -130 96 -129
rect 96 -130 97 -129
rect 97 -130 98 -129
rect 98 -130 99 -129
rect 99 -130 100 -129
rect 100 -130 101 -129
rect 101 -130 102 -129
rect 102 -130 103 -129
rect 103 -130 104 -129
rect 104 -130 105 -129
rect 105 -130 106 -129
rect 106 -130 107 -129
rect 107 -130 108 -129
rect 108 -130 109 -129
rect 109 -130 110 -129
rect 110 -130 111 -129
rect 111 -130 112 -129
rect 112 -130 113 -129
rect 113 -130 114 -129
rect 114 -130 115 -129
rect 115 -130 116 -129
rect 116 -130 117 -129
rect 117 -130 118 -129
rect 118 -130 119 -129
rect 119 -130 120 -129
rect 120 -130 121 -129
rect 121 -130 122 -129
rect 122 -130 123 -129
rect 123 -130 124 -129
rect 124 -130 125 -129
rect 125 -130 126 -129
rect 126 -130 127 -129
rect 127 -130 128 -129
rect 128 -130 129 -129
rect 129 -130 130 -129
rect 130 -130 131 -129
rect 131 -130 132 -129
rect 132 -130 133 -129
rect 133 -130 134 -129
rect 134 -130 135 -129
rect 135 -130 136 -129
rect 136 -130 137 -129
rect 137 -130 138 -129
rect 138 -130 139 -129
rect 139 -130 140 -129
rect 140 -130 141 -129
rect 141 -130 142 -129
rect 142 -130 143 -129
rect 143 -130 144 -129
rect 144 -130 145 -129
rect 145 -130 146 -129
rect 146 -130 147 -129
rect 147 -130 148 -129
rect 148 -130 149 -129
rect 149 -130 150 -129
rect 150 -130 151 -129
rect 151 -130 152 -129
rect 152 -130 153 -129
rect 153 -130 154 -129
rect 154 -130 155 -129
rect 155 -130 156 -129
rect 156 -130 157 -129
rect 157 -130 158 -129
rect 158 -130 159 -129
rect 159 -130 160 -129
rect 160 -130 161 -129
rect 161 -130 162 -129
rect 162 -130 163 -129
rect 163 -130 164 -129
rect 164 -130 165 -129
rect 165 -130 166 -129
rect 166 -130 167 -129
rect 167 -130 168 -129
rect 168 -130 169 -129
rect 169 -130 170 -129
rect 170 -130 171 -129
rect 171 -130 172 -129
rect 172 -130 173 -129
rect 173 -130 174 -129
rect 174 -130 175 -129
rect 175 -130 176 -129
rect 176 -130 177 -129
rect 177 -130 178 -129
rect 178 -130 179 -129
rect 179 -130 180 -129
rect 180 -130 181 -129
rect 181 -130 182 -129
rect 182 -130 183 -129
rect 183 -130 184 -129
rect 184 -130 185 -129
rect 185 -130 186 -129
rect 186 -130 187 -129
rect 187 -130 188 -129
rect 188 -130 189 -129
rect 189 -130 190 -129
rect 190 -130 191 -129
rect 191 -130 192 -129
rect 192 -130 193 -129
rect 193 -130 194 -129
rect 194 -130 195 -129
rect 195 -130 196 -129
rect 196 -130 197 -129
rect 197 -130 198 -129
rect 198 -130 199 -129
rect 199 -130 200 -129
rect 200 -130 201 -129
rect 201 -130 202 -129
rect 202 -130 203 -129
rect 203 -130 204 -129
rect 204 -130 205 -129
rect 205 -130 206 -129
rect 206 -130 207 -129
rect 207 -130 208 -129
rect 208 -130 209 -129
rect 209 -130 210 -129
rect 210 -130 211 -129
rect 211 -130 212 -129
rect 212 -130 213 -129
rect 213 -130 214 -129
rect 214 -130 215 -129
rect 215 -130 216 -129
rect 216 -130 217 -129
rect 217 -130 218 -129
rect 218 -130 219 -129
rect 219 -130 220 -129
rect 220 -130 221 -129
rect 221 -130 222 -129
rect 222 -130 223 -129
rect 223 -130 224 -129
rect 224 -130 225 -129
rect 225 -130 226 -129
rect 226 -130 227 -129
rect 227 -130 228 -129
rect 228 -130 229 -129
rect 229 -130 230 -129
rect 230 -130 231 -129
rect 231 -130 232 -129
rect 232 -130 233 -129
rect 233 -130 234 -129
rect 234 -130 235 -129
rect 235 -130 236 -129
rect 236 -130 237 -129
rect 237 -130 238 -129
rect 238 -130 239 -129
rect 239 -130 240 -129
rect 240 -130 241 -129
rect 241 -130 242 -129
rect 242 -130 243 -129
rect 243 -130 244 -129
rect 244 -130 245 -129
rect 245 -130 246 -129
rect 246 -130 247 -129
rect 247 -130 248 -129
rect 248 -130 249 -129
rect 249 -130 250 -129
rect 250 -130 251 -129
rect 251 -130 252 -129
rect 252 -130 253 -129
rect 253 -130 254 -129
rect 254 -130 255 -129
rect 255 -130 256 -129
rect 256 -130 257 -129
rect 257 -130 258 -129
rect 258 -130 259 -129
rect 259 -130 260 -129
rect 260 -130 261 -129
rect 261 -130 262 -129
rect 262 -130 263 -129
rect 263 -130 264 -129
rect 264 -130 265 -129
rect 265 -130 266 -129
rect 266 -130 267 -129
rect 267 -130 268 -129
rect 268 -130 269 -129
rect 269 -130 270 -129
rect 270 -130 271 -129
rect 271 -130 272 -129
rect 272 -130 273 -129
rect 273 -130 274 -129
rect 274 -130 275 -129
rect 275 -130 276 -129
rect 276 -130 277 -129
rect 277 -130 278 -129
rect 278 -130 279 -129
rect 279 -130 280 -129
rect 280 -130 281 -129
rect 281 -130 282 -129
rect 282 -130 283 -129
rect 283 -130 284 -129
rect 284 -130 285 -129
rect 285 -130 286 -129
rect 286 -130 287 -129
rect 287 -130 288 -129
rect 288 -130 289 -129
rect 289 -130 290 -129
rect 290 -130 291 -129
rect 291 -130 292 -129
rect 292 -130 293 -129
rect 293 -130 294 -129
rect 294 -130 295 -129
rect 295 -130 296 -129
rect 296 -130 297 -129
rect 297 -130 298 -129
rect 298 -130 299 -129
rect 299 -130 300 -129
rect 300 -130 301 -129
rect 301 -130 302 -129
rect 302 -130 303 -129
rect 303 -130 304 -129
rect 304 -130 305 -129
rect 305 -130 306 -129
rect 306 -130 307 -129
rect 307 -130 308 -129
rect 308 -130 309 -129
rect 309 -130 310 -129
rect 310 -130 311 -129
rect 311 -130 312 -129
rect 312 -130 313 -129
rect 313 -130 314 -129
rect 314 -130 315 -129
rect 315 -130 316 -129
rect 316 -130 317 -129
rect 317 -130 318 -129
rect 318 -130 319 -129
rect 319 -130 320 -129
rect 320 -130 321 -129
rect 321 -130 322 -129
rect 322 -130 323 -129
rect 323 -130 324 -129
rect 324 -130 325 -129
rect 325 -130 326 -129
rect 326 -130 327 -129
rect 327 -130 328 -129
rect 328 -130 329 -129
rect 329 -130 330 -129
rect 330 -130 331 -129
rect 331 -130 332 -129
rect 332 -130 333 -129
rect 333 -130 334 -129
rect 334 -130 335 -129
rect 335 -130 336 -129
rect 336 -130 337 -129
rect 337 -130 338 -129
rect 338 -130 339 -129
rect 339 -130 340 -129
rect 340 -130 341 -129
rect 341 -130 342 -129
rect 342 -130 343 -129
rect 343 -130 344 -129
rect 344 -130 345 -129
rect 345 -130 346 -129
rect 346 -130 347 -129
rect 347 -130 348 -129
rect 348 -130 349 -129
rect 349 -130 350 -129
rect 350 -130 351 -129
rect 351 -130 352 -129
rect 352 -130 353 -129
rect 353 -130 354 -129
rect 354 -130 355 -129
rect 355 -130 356 -129
rect 356 -130 357 -129
rect 357 -130 358 -129
rect 358 -130 359 -129
rect 359 -130 360 -129
rect 360 -130 361 -129
rect 361 -130 362 -129
rect 362 -130 363 -129
rect 363 -130 364 -129
rect 364 -130 365 -129
rect 365 -130 366 -129
rect 366 -130 367 -129
rect 367 -130 368 -129
rect 368 -130 369 -129
rect 369 -130 370 -129
rect 370 -130 371 -129
rect 371 -130 372 -129
rect 372 -130 373 -129
rect 373 -130 374 -129
rect 374 -130 375 -129
rect 375 -130 376 -129
rect 376 -130 377 -129
rect 377 -130 378 -129
rect 378 -130 379 -129
rect 379 -130 380 -129
rect 380 -130 381 -129
rect 381 -130 382 -129
rect 382 -130 383 -129
rect 383 -130 384 -129
rect 384 -130 385 -129
rect 385 -130 386 -129
rect 386 -130 387 -129
rect 387 -130 388 -129
rect 388 -130 389 -129
rect 389 -130 390 -129
rect 390 -130 391 -129
rect 391 -130 392 -129
rect 392 -130 393 -129
rect 393 -130 394 -129
rect 394 -130 395 -129
rect 395 -130 396 -129
rect 396 -130 397 -129
rect 397 -130 398 -129
rect 398 -130 399 -129
rect 399 -130 400 -129
rect 400 -130 401 -129
rect 401 -130 402 -129
rect 402 -130 403 -129
rect 403 -130 404 -129
rect 404 -130 405 -129
rect 405 -130 406 -129
rect 406 -130 407 -129
rect 407 -130 408 -129
rect 408 -130 409 -129
rect 409 -130 410 -129
rect 410 -130 411 -129
rect 411 -130 412 -129
rect 412 -130 413 -129
rect 413 -130 414 -129
rect 414 -130 415 -129
rect 415 -130 416 -129
rect 416 -130 417 -129
rect 417 -130 418 -129
rect 418 -130 419 -129
rect 419 -130 420 -129
rect 420 -130 421 -129
rect 421 -130 422 -129
rect 422 -130 423 -129
rect 423 -130 424 -129
rect 424 -130 425 -129
rect 425 -130 426 -129
rect 426 -130 427 -129
rect 427 -130 428 -129
rect 428 -130 429 -129
rect 429 -130 430 -129
rect 430 -130 431 -129
rect 431 -130 432 -129
rect 432 -130 433 -129
rect 433 -130 434 -129
rect 434 -130 435 -129
rect 435 -130 436 -129
rect 436 -130 437 -129
rect 437 -130 438 -129
rect 438 -130 439 -129
rect 439 -130 440 -129
rect 440 -130 441 -129
rect 441 -130 442 -129
rect 442 -130 443 -129
rect 443 -130 444 -129
rect 444 -130 445 -129
rect 445 -130 446 -129
rect 446 -130 447 -129
rect 447 -130 448 -129
rect 448 -130 449 -129
rect 449 -130 450 -129
rect 450 -130 451 -129
rect 451 -130 452 -129
rect 452 -130 453 -129
rect 453 -130 454 -129
rect 454 -130 455 -129
rect 455 -130 456 -129
rect 456 -130 457 -129
rect 457 -130 458 -129
rect 458 -130 459 -129
rect 459 -130 460 -129
rect 460 -130 461 -129
rect 461 -130 462 -129
rect 462 -130 463 -129
rect 463 -130 464 -129
rect 464 -130 465 -129
rect 465 -130 466 -129
rect 466 -130 467 -129
rect 467 -130 468 -129
rect 468 -130 469 -129
rect 469 -130 470 -129
rect 470 -130 471 -129
rect 471 -130 472 -129
rect 472 -130 473 -129
rect 473 -130 474 -129
rect 474 -130 475 -129
rect 475 -130 476 -129
rect 476 -130 477 -129
rect 477 -130 478 -129
rect 478 -130 479 -129
rect 479 -130 480 -129
rect 2 -131 3 -130
rect 3 -131 4 -130
rect 4 -131 5 -130
rect 5 -131 6 -130
rect 6 -131 7 -130
rect 7 -131 8 -130
rect 8 -131 9 -130
rect 9 -131 10 -130
rect 10 -131 11 -130
rect 11 -131 12 -130
rect 12 -131 13 -130
rect 13 -131 14 -130
rect 14 -131 15 -130
rect 15 -131 16 -130
rect 16 -131 17 -130
rect 17 -131 18 -130
rect 18 -131 19 -130
rect 19 -131 20 -130
rect 20 -131 21 -130
rect 21 -131 22 -130
rect 22 -131 23 -130
rect 23 -131 24 -130
rect 24 -131 25 -130
rect 25 -131 26 -130
rect 26 -131 27 -130
rect 27 -131 28 -130
rect 28 -131 29 -130
rect 29 -131 30 -130
rect 30 -131 31 -130
rect 31 -131 32 -130
rect 32 -131 33 -130
rect 33 -131 34 -130
rect 34 -131 35 -130
rect 35 -131 36 -130
rect 36 -131 37 -130
rect 37 -131 38 -130
rect 38 -131 39 -130
rect 39 -131 40 -130
rect 40 -131 41 -130
rect 41 -131 42 -130
rect 42 -131 43 -130
rect 43 -131 44 -130
rect 44 -131 45 -130
rect 45 -131 46 -130
rect 46 -131 47 -130
rect 47 -131 48 -130
rect 48 -131 49 -130
rect 49 -131 50 -130
rect 50 -131 51 -130
rect 51 -131 52 -130
rect 52 -131 53 -130
rect 53 -131 54 -130
rect 54 -131 55 -130
rect 55 -131 56 -130
rect 56 -131 57 -130
rect 57 -131 58 -130
rect 58 -131 59 -130
rect 59 -131 60 -130
rect 60 -131 61 -130
rect 61 -131 62 -130
rect 62 -131 63 -130
rect 63 -131 64 -130
rect 64 -131 65 -130
rect 65 -131 66 -130
rect 66 -131 67 -130
rect 67 -131 68 -130
rect 68 -131 69 -130
rect 69 -131 70 -130
rect 70 -131 71 -130
rect 71 -131 72 -130
rect 72 -131 73 -130
rect 73 -131 74 -130
rect 74 -131 75 -130
rect 75 -131 76 -130
rect 76 -131 77 -130
rect 77 -131 78 -130
rect 78 -131 79 -130
rect 79 -131 80 -130
rect 80 -131 81 -130
rect 81 -131 82 -130
rect 82 -131 83 -130
rect 83 -131 84 -130
rect 84 -131 85 -130
rect 85 -131 86 -130
rect 86 -131 87 -130
rect 87 -131 88 -130
rect 88 -131 89 -130
rect 89 -131 90 -130
rect 90 -131 91 -130
rect 91 -131 92 -130
rect 92 -131 93 -130
rect 93 -131 94 -130
rect 94 -131 95 -130
rect 95 -131 96 -130
rect 96 -131 97 -130
rect 97 -131 98 -130
rect 98 -131 99 -130
rect 99 -131 100 -130
rect 100 -131 101 -130
rect 101 -131 102 -130
rect 102 -131 103 -130
rect 103 -131 104 -130
rect 104 -131 105 -130
rect 105 -131 106 -130
rect 106 -131 107 -130
rect 107 -131 108 -130
rect 108 -131 109 -130
rect 109 -131 110 -130
rect 110 -131 111 -130
rect 111 -131 112 -130
rect 112 -131 113 -130
rect 113 -131 114 -130
rect 114 -131 115 -130
rect 115 -131 116 -130
rect 116 -131 117 -130
rect 117 -131 118 -130
rect 118 -131 119 -130
rect 119 -131 120 -130
rect 120 -131 121 -130
rect 121 -131 122 -130
rect 122 -131 123 -130
rect 123 -131 124 -130
rect 124 -131 125 -130
rect 125 -131 126 -130
rect 126 -131 127 -130
rect 127 -131 128 -130
rect 128 -131 129 -130
rect 129 -131 130 -130
rect 130 -131 131 -130
rect 131 -131 132 -130
rect 132 -131 133 -130
rect 133 -131 134 -130
rect 134 -131 135 -130
rect 135 -131 136 -130
rect 136 -131 137 -130
rect 137 -131 138 -130
rect 138 -131 139 -130
rect 139 -131 140 -130
rect 140 -131 141 -130
rect 141 -131 142 -130
rect 142 -131 143 -130
rect 143 -131 144 -130
rect 144 -131 145 -130
rect 145 -131 146 -130
rect 146 -131 147 -130
rect 147 -131 148 -130
rect 148 -131 149 -130
rect 149 -131 150 -130
rect 150 -131 151 -130
rect 151 -131 152 -130
rect 152 -131 153 -130
rect 153 -131 154 -130
rect 154 -131 155 -130
rect 155 -131 156 -130
rect 156 -131 157 -130
rect 157 -131 158 -130
rect 158 -131 159 -130
rect 159 -131 160 -130
rect 160 -131 161 -130
rect 161 -131 162 -130
rect 162 -131 163 -130
rect 163 -131 164 -130
rect 164 -131 165 -130
rect 165 -131 166 -130
rect 166 -131 167 -130
rect 167 -131 168 -130
rect 168 -131 169 -130
rect 169 -131 170 -130
rect 170 -131 171 -130
rect 171 -131 172 -130
rect 172 -131 173 -130
rect 173 -131 174 -130
rect 174 -131 175 -130
rect 175 -131 176 -130
rect 176 -131 177 -130
rect 177 -131 178 -130
rect 178 -131 179 -130
rect 179 -131 180 -130
rect 180 -131 181 -130
rect 181 -131 182 -130
rect 182 -131 183 -130
rect 183 -131 184 -130
rect 184 -131 185 -130
rect 185 -131 186 -130
rect 186 -131 187 -130
rect 187 -131 188 -130
rect 188 -131 189 -130
rect 189 -131 190 -130
rect 190 -131 191 -130
rect 191 -131 192 -130
rect 192 -131 193 -130
rect 193 -131 194 -130
rect 194 -131 195 -130
rect 195 -131 196 -130
rect 196 -131 197 -130
rect 197 -131 198 -130
rect 198 -131 199 -130
rect 199 -131 200 -130
rect 200 -131 201 -130
rect 201 -131 202 -130
rect 202 -131 203 -130
rect 203 -131 204 -130
rect 204 -131 205 -130
rect 205 -131 206 -130
rect 206 -131 207 -130
rect 207 -131 208 -130
rect 208 -131 209 -130
rect 209 -131 210 -130
rect 210 -131 211 -130
rect 211 -131 212 -130
rect 212 -131 213 -130
rect 213 -131 214 -130
rect 214 -131 215 -130
rect 215 -131 216 -130
rect 216 -131 217 -130
rect 217 -131 218 -130
rect 218 -131 219 -130
rect 219 -131 220 -130
rect 220 -131 221 -130
rect 221 -131 222 -130
rect 222 -131 223 -130
rect 223 -131 224 -130
rect 224 -131 225 -130
rect 225 -131 226 -130
rect 226 -131 227 -130
rect 227 -131 228 -130
rect 228 -131 229 -130
rect 229 -131 230 -130
rect 230 -131 231 -130
rect 231 -131 232 -130
rect 232 -131 233 -130
rect 233 -131 234 -130
rect 234 -131 235 -130
rect 235 -131 236 -130
rect 236 -131 237 -130
rect 237 -131 238 -130
rect 238 -131 239 -130
rect 239 -131 240 -130
rect 240 -131 241 -130
rect 241 -131 242 -130
rect 242 -131 243 -130
rect 243 -131 244 -130
rect 244 -131 245 -130
rect 245 -131 246 -130
rect 246 -131 247 -130
rect 247 -131 248 -130
rect 248 -131 249 -130
rect 249 -131 250 -130
rect 250 -131 251 -130
rect 251 -131 252 -130
rect 252 -131 253 -130
rect 253 -131 254 -130
rect 254 -131 255 -130
rect 255 -131 256 -130
rect 256 -131 257 -130
rect 257 -131 258 -130
rect 258 -131 259 -130
rect 259 -131 260 -130
rect 260 -131 261 -130
rect 261 -131 262 -130
rect 262 -131 263 -130
rect 263 -131 264 -130
rect 264 -131 265 -130
rect 265 -131 266 -130
rect 266 -131 267 -130
rect 267 -131 268 -130
rect 268 -131 269 -130
rect 269 -131 270 -130
rect 270 -131 271 -130
rect 271 -131 272 -130
rect 272 -131 273 -130
rect 273 -131 274 -130
rect 274 -131 275 -130
rect 275 -131 276 -130
rect 276 -131 277 -130
rect 277 -131 278 -130
rect 278 -131 279 -130
rect 279 -131 280 -130
rect 280 -131 281 -130
rect 281 -131 282 -130
rect 282 -131 283 -130
rect 283 -131 284 -130
rect 284 -131 285 -130
rect 285 -131 286 -130
rect 286 -131 287 -130
rect 287 -131 288 -130
rect 288 -131 289 -130
rect 289 -131 290 -130
rect 290 -131 291 -130
rect 291 -131 292 -130
rect 292 -131 293 -130
rect 293 -131 294 -130
rect 294 -131 295 -130
rect 295 -131 296 -130
rect 296 -131 297 -130
rect 297 -131 298 -130
rect 298 -131 299 -130
rect 299 -131 300 -130
rect 300 -131 301 -130
rect 301 -131 302 -130
rect 302 -131 303 -130
rect 303 -131 304 -130
rect 304 -131 305 -130
rect 305 -131 306 -130
rect 306 -131 307 -130
rect 307 -131 308 -130
rect 308 -131 309 -130
rect 309 -131 310 -130
rect 310 -131 311 -130
rect 311 -131 312 -130
rect 312 -131 313 -130
rect 313 -131 314 -130
rect 314 -131 315 -130
rect 315 -131 316 -130
rect 316 -131 317 -130
rect 317 -131 318 -130
rect 318 -131 319 -130
rect 319 -131 320 -130
rect 320 -131 321 -130
rect 321 -131 322 -130
rect 322 -131 323 -130
rect 323 -131 324 -130
rect 324 -131 325 -130
rect 325 -131 326 -130
rect 326 -131 327 -130
rect 327 -131 328 -130
rect 328 -131 329 -130
rect 329 -131 330 -130
rect 330 -131 331 -130
rect 331 -131 332 -130
rect 332 -131 333 -130
rect 333 -131 334 -130
rect 334 -131 335 -130
rect 335 -131 336 -130
rect 336 -131 337 -130
rect 337 -131 338 -130
rect 338 -131 339 -130
rect 339 -131 340 -130
rect 340 -131 341 -130
rect 341 -131 342 -130
rect 342 -131 343 -130
rect 343 -131 344 -130
rect 344 -131 345 -130
rect 345 -131 346 -130
rect 346 -131 347 -130
rect 347 -131 348 -130
rect 348 -131 349 -130
rect 349 -131 350 -130
rect 350 -131 351 -130
rect 351 -131 352 -130
rect 352 -131 353 -130
rect 353 -131 354 -130
rect 354 -131 355 -130
rect 355 -131 356 -130
rect 356 -131 357 -130
rect 357 -131 358 -130
rect 358 -131 359 -130
rect 359 -131 360 -130
rect 360 -131 361 -130
rect 361 -131 362 -130
rect 362 -131 363 -130
rect 363 -131 364 -130
rect 364 -131 365 -130
rect 365 -131 366 -130
rect 366 -131 367 -130
rect 367 -131 368 -130
rect 368 -131 369 -130
rect 369 -131 370 -130
rect 370 -131 371 -130
rect 371 -131 372 -130
rect 372 -131 373 -130
rect 373 -131 374 -130
rect 374 -131 375 -130
rect 375 -131 376 -130
rect 376 -131 377 -130
rect 377 -131 378 -130
rect 378 -131 379 -130
rect 379 -131 380 -130
rect 380 -131 381 -130
rect 381 -131 382 -130
rect 382 -131 383 -130
rect 383 -131 384 -130
rect 384 -131 385 -130
rect 385 -131 386 -130
rect 386 -131 387 -130
rect 387 -131 388 -130
rect 388 -131 389 -130
rect 389 -131 390 -130
rect 390 -131 391 -130
rect 391 -131 392 -130
rect 392 -131 393 -130
rect 393 -131 394 -130
rect 394 -131 395 -130
rect 395 -131 396 -130
rect 396 -131 397 -130
rect 397 -131 398 -130
rect 398 -131 399 -130
rect 399 -131 400 -130
rect 400 -131 401 -130
rect 401 -131 402 -130
rect 402 -131 403 -130
rect 403 -131 404 -130
rect 404 -131 405 -130
rect 405 -131 406 -130
rect 406 -131 407 -130
rect 407 -131 408 -130
rect 408 -131 409 -130
rect 409 -131 410 -130
rect 410 -131 411 -130
rect 411 -131 412 -130
rect 412 -131 413 -130
rect 413 -131 414 -130
rect 414 -131 415 -130
rect 415 -131 416 -130
rect 416 -131 417 -130
rect 417 -131 418 -130
rect 418 -131 419 -130
rect 419 -131 420 -130
rect 420 -131 421 -130
rect 421 -131 422 -130
rect 422 -131 423 -130
rect 423 -131 424 -130
rect 424 -131 425 -130
rect 425 -131 426 -130
rect 426 -131 427 -130
rect 427 -131 428 -130
rect 428 -131 429 -130
rect 429 -131 430 -130
rect 430 -131 431 -130
rect 431 -131 432 -130
rect 432 -131 433 -130
rect 433 -131 434 -130
rect 434 -131 435 -130
rect 435 -131 436 -130
rect 436 -131 437 -130
rect 437 -131 438 -130
rect 438 -131 439 -130
rect 439 -131 440 -130
rect 440 -131 441 -130
rect 441 -131 442 -130
rect 442 -131 443 -130
rect 443 -131 444 -130
rect 444 -131 445 -130
rect 445 -131 446 -130
rect 446 -131 447 -130
rect 447 -131 448 -130
rect 448 -131 449 -130
rect 449 -131 450 -130
rect 450 -131 451 -130
rect 451 -131 452 -130
rect 452 -131 453 -130
rect 453 -131 454 -130
rect 454 -131 455 -130
rect 455 -131 456 -130
rect 456 -131 457 -130
rect 457 -131 458 -130
rect 458 -131 459 -130
rect 459 -131 460 -130
rect 460 -131 461 -130
rect 461 -131 462 -130
rect 462 -131 463 -130
rect 463 -131 464 -130
rect 464 -131 465 -130
rect 465 -131 466 -130
rect 466 -131 467 -130
rect 467 -131 468 -130
rect 468 -131 469 -130
rect 469 -131 470 -130
rect 470 -131 471 -130
rect 471 -131 472 -130
rect 472 -131 473 -130
rect 473 -131 474 -130
rect 474 -131 475 -130
rect 475 -131 476 -130
rect 476 -131 477 -130
rect 477 -131 478 -130
rect 478 -131 479 -130
rect 479 -131 480 -130
rect 2 -132 3 -131
rect 3 -132 4 -131
rect 4 -132 5 -131
rect 5 -132 6 -131
rect 6 -132 7 -131
rect 7 -132 8 -131
rect 8 -132 9 -131
rect 9 -132 10 -131
rect 10 -132 11 -131
rect 11 -132 12 -131
rect 12 -132 13 -131
rect 13 -132 14 -131
rect 14 -132 15 -131
rect 15 -132 16 -131
rect 16 -132 17 -131
rect 17 -132 18 -131
rect 18 -132 19 -131
rect 19 -132 20 -131
rect 20 -132 21 -131
rect 21 -132 22 -131
rect 22 -132 23 -131
rect 23 -132 24 -131
rect 24 -132 25 -131
rect 25 -132 26 -131
rect 26 -132 27 -131
rect 27 -132 28 -131
rect 28 -132 29 -131
rect 29 -132 30 -131
rect 30 -132 31 -131
rect 31 -132 32 -131
rect 32 -132 33 -131
rect 33 -132 34 -131
rect 34 -132 35 -131
rect 35 -132 36 -131
rect 36 -132 37 -131
rect 37 -132 38 -131
rect 38 -132 39 -131
rect 39 -132 40 -131
rect 40 -132 41 -131
rect 41 -132 42 -131
rect 42 -132 43 -131
rect 43 -132 44 -131
rect 44 -132 45 -131
rect 45 -132 46 -131
rect 46 -132 47 -131
rect 47 -132 48 -131
rect 48 -132 49 -131
rect 49 -132 50 -131
rect 50 -132 51 -131
rect 51 -132 52 -131
rect 52 -132 53 -131
rect 53 -132 54 -131
rect 54 -132 55 -131
rect 55 -132 56 -131
rect 56 -132 57 -131
rect 57 -132 58 -131
rect 58 -132 59 -131
rect 59 -132 60 -131
rect 60 -132 61 -131
rect 61 -132 62 -131
rect 62 -132 63 -131
rect 63 -132 64 -131
rect 64 -132 65 -131
rect 65 -132 66 -131
rect 66 -132 67 -131
rect 67 -132 68 -131
rect 68 -132 69 -131
rect 69 -132 70 -131
rect 70 -132 71 -131
rect 71 -132 72 -131
rect 72 -132 73 -131
rect 73 -132 74 -131
rect 74 -132 75 -131
rect 75 -132 76 -131
rect 76 -132 77 -131
rect 77 -132 78 -131
rect 78 -132 79 -131
rect 79 -132 80 -131
rect 80 -132 81 -131
rect 81 -132 82 -131
rect 82 -132 83 -131
rect 83 -132 84 -131
rect 84 -132 85 -131
rect 85 -132 86 -131
rect 86 -132 87 -131
rect 87 -132 88 -131
rect 88 -132 89 -131
rect 89 -132 90 -131
rect 90 -132 91 -131
rect 91 -132 92 -131
rect 92 -132 93 -131
rect 93 -132 94 -131
rect 94 -132 95 -131
rect 95 -132 96 -131
rect 96 -132 97 -131
rect 97 -132 98 -131
rect 98 -132 99 -131
rect 99 -132 100 -131
rect 100 -132 101 -131
rect 101 -132 102 -131
rect 102 -132 103 -131
rect 103 -132 104 -131
rect 104 -132 105 -131
rect 105 -132 106 -131
rect 106 -132 107 -131
rect 107 -132 108 -131
rect 108 -132 109 -131
rect 109 -132 110 -131
rect 110 -132 111 -131
rect 111 -132 112 -131
rect 112 -132 113 -131
rect 113 -132 114 -131
rect 114 -132 115 -131
rect 115 -132 116 -131
rect 116 -132 117 -131
rect 117 -132 118 -131
rect 118 -132 119 -131
rect 119 -132 120 -131
rect 120 -132 121 -131
rect 121 -132 122 -131
rect 122 -132 123 -131
rect 123 -132 124 -131
rect 124 -132 125 -131
rect 125 -132 126 -131
rect 126 -132 127 -131
rect 127 -132 128 -131
rect 128 -132 129 -131
rect 129 -132 130 -131
rect 130 -132 131 -131
rect 131 -132 132 -131
rect 132 -132 133 -131
rect 133 -132 134 -131
rect 134 -132 135 -131
rect 135 -132 136 -131
rect 136 -132 137 -131
rect 137 -132 138 -131
rect 138 -132 139 -131
rect 139 -132 140 -131
rect 140 -132 141 -131
rect 141 -132 142 -131
rect 142 -132 143 -131
rect 143 -132 144 -131
rect 144 -132 145 -131
rect 145 -132 146 -131
rect 146 -132 147 -131
rect 147 -132 148 -131
rect 148 -132 149 -131
rect 149 -132 150 -131
rect 150 -132 151 -131
rect 151 -132 152 -131
rect 152 -132 153 -131
rect 153 -132 154 -131
rect 154 -132 155 -131
rect 155 -132 156 -131
rect 156 -132 157 -131
rect 157 -132 158 -131
rect 158 -132 159 -131
rect 159 -132 160 -131
rect 160 -132 161 -131
rect 161 -132 162 -131
rect 162 -132 163 -131
rect 163 -132 164 -131
rect 164 -132 165 -131
rect 165 -132 166 -131
rect 166 -132 167 -131
rect 167 -132 168 -131
rect 168 -132 169 -131
rect 169 -132 170 -131
rect 170 -132 171 -131
rect 171 -132 172 -131
rect 172 -132 173 -131
rect 173 -132 174 -131
rect 174 -132 175 -131
rect 175 -132 176 -131
rect 176 -132 177 -131
rect 177 -132 178 -131
rect 178 -132 179 -131
rect 179 -132 180 -131
rect 180 -132 181 -131
rect 181 -132 182 -131
rect 182 -132 183 -131
rect 183 -132 184 -131
rect 184 -132 185 -131
rect 185 -132 186 -131
rect 186 -132 187 -131
rect 187 -132 188 -131
rect 188 -132 189 -131
rect 189 -132 190 -131
rect 190 -132 191 -131
rect 191 -132 192 -131
rect 192 -132 193 -131
rect 193 -132 194 -131
rect 194 -132 195 -131
rect 195 -132 196 -131
rect 196 -132 197 -131
rect 197 -132 198 -131
rect 198 -132 199 -131
rect 199 -132 200 -131
rect 200 -132 201 -131
rect 201 -132 202 -131
rect 202 -132 203 -131
rect 203 -132 204 -131
rect 204 -132 205 -131
rect 205 -132 206 -131
rect 206 -132 207 -131
rect 207 -132 208 -131
rect 208 -132 209 -131
rect 209 -132 210 -131
rect 210 -132 211 -131
rect 211 -132 212 -131
rect 212 -132 213 -131
rect 213 -132 214 -131
rect 214 -132 215 -131
rect 215 -132 216 -131
rect 216 -132 217 -131
rect 217 -132 218 -131
rect 218 -132 219 -131
rect 219 -132 220 -131
rect 220 -132 221 -131
rect 221 -132 222 -131
rect 222 -132 223 -131
rect 223 -132 224 -131
rect 224 -132 225 -131
rect 225 -132 226 -131
rect 226 -132 227 -131
rect 227 -132 228 -131
rect 228 -132 229 -131
rect 229 -132 230 -131
rect 230 -132 231 -131
rect 231 -132 232 -131
rect 232 -132 233 -131
rect 233 -132 234 -131
rect 234 -132 235 -131
rect 235 -132 236 -131
rect 236 -132 237 -131
rect 237 -132 238 -131
rect 238 -132 239 -131
rect 239 -132 240 -131
rect 240 -132 241 -131
rect 241 -132 242 -131
rect 242 -132 243 -131
rect 243 -132 244 -131
rect 244 -132 245 -131
rect 245 -132 246 -131
rect 246 -132 247 -131
rect 247 -132 248 -131
rect 248 -132 249 -131
rect 249 -132 250 -131
rect 250 -132 251 -131
rect 251 -132 252 -131
rect 252 -132 253 -131
rect 253 -132 254 -131
rect 254 -132 255 -131
rect 255 -132 256 -131
rect 256 -132 257 -131
rect 257 -132 258 -131
rect 258 -132 259 -131
rect 259 -132 260 -131
rect 260 -132 261 -131
rect 261 -132 262 -131
rect 262 -132 263 -131
rect 263 -132 264 -131
rect 264 -132 265 -131
rect 265 -132 266 -131
rect 266 -132 267 -131
rect 267 -132 268 -131
rect 268 -132 269 -131
rect 269 -132 270 -131
rect 270 -132 271 -131
rect 271 -132 272 -131
rect 272 -132 273 -131
rect 273 -132 274 -131
rect 274 -132 275 -131
rect 275 -132 276 -131
rect 276 -132 277 -131
rect 277 -132 278 -131
rect 278 -132 279 -131
rect 279 -132 280 -131
rect 280 -132 281 -131
rect 281 -132 282 -131
rect 282 -132 283 -131
rect 283 -132 284 -131
rect 284 -132 285 -131
rect 285 -132 286 -131
rect 286 -132 287 -131
rect 287 -132 288 -131
rect 288 -132 289 -131
rect 289 -132 290 -131
rect 290 -132 291 -131
rect 291 -132 292 -131
rect 292 -132 293 -131
rect 293 -132 294 -131
rect 294 -132 295 -131
rect 295 -132 296 -131
rect 296 -132 297 -131
rect 297 -132 298 -131
rect 298 -132 299 -131
rect 299 -132 300 -131
rect 300 -132 301 -131
rect 301 -132 302 -131
rect 302 -132 303 -131
rect 303 -132 304 -131
rect 304 -132 305 -131
rect 305 -132 306 -131
rect 306 -132 307 -131
rect 307 -132 308 -131
rect 308 -132 309 -131
rect 309 -132 310 -131
rect 310 -132 311 -131
rect 311 -132 312 -131
rect 312 -132 313 -131
rect 313 -132 314 -131
rect 314 -132 315 -131
rect 315 -132 316 -131
rect 316 -132 317 -131
rect 317 -132 318 -131
rect 318 -132 319 -131
rect 319 -132 320 -131
rect 320 -132 321 -131
rect 321 -132 322 -131
rect 322 -132 323 -131
rect 323 -132 324 -131
rect 324 -132 325 -131
rect 325 -132 326 -131
rect 326 -132 327 -131
rect 327 -132 328 -131
rect 328 -132 329 -131
rect 329 -132 330 -131
rect 330 -132 331 -131
rect 331 -132 332 -131
rect 332 -132 333 -131
rect 333 -132 334 -131
rect 334 -132 335 -131
rect 335 -132 336 -131
rect 336 -132 337 -131
rect 337 -132 338 -131
rect 338 -132 339 -131
rect 339 -132 340 -131
rect 340 -132 341 -131
rect 341 -132 342 -131
rect 342 -132 343 -131
rect 343 -132 344 -131
rect 344 -132 345 -131
rect 345 -132 346 -131
rect 346 -132 347 -131
rect 347 -132 348 -131
rect 348 -132 349 -131
rect 349 -132 350 -131
rect 350 -132 351 -131
rect 351 -132 352 -131
rect 352 -132 353 -131
rect 353 -132 354 -131
rect 354 -132 355 -131
rect 355 -132 356 -131
rect 356 -132 357 -131
rect 357 -132 358 -131
rect 358 -132 359 -131
rect 359 -132 360 -131
rect 360 -132 361 -131
rect 361 -132 362 -131
rect 362 -132 363 -131
rect 363 -132 364 -131
rect 364 -132 365 -131
rect 365 -132 366 -131
rect 366 -132 367 -131
rect 367 -132 368 -131
rect 368 -132 369 -131
rect 369 -132 370 -131
rect 370 -132 371 -131
rect 371 -132 372 -131
rect 372 -132 373 -131
rect 373 -132 374 -131
rect 374 -132 375 -131
rect 375 -132 376 -131
rect 376 -132 377 -131
rect 377 -132 378 -131
rect 378 -132 379 -131
rect 379 -132 380 -131
rect 380 -132 381 -131
rect 381 -132 382 -131
rect 382 -132 383 -131
rect 383 -132 384 -131
rect 384 -132 385 -131
rect 385 -132 386 -131
rect 386 -132 387 -131
rect 387 -132 388 -131
rect 388 -132 389 -131
rect 389 -132 390 -131
rect 390 -132 391 -131
rect 391 -132 392 -131
rect 392 -132 393 -131
rect 393 -132 394 -131
rect 394 -132 395 -131
rect 395 -132 396 -131
rect 396 -132 397 -131
rect 397 -132 398 -131
rect 398 -132 399 -131
rect 399 -132 400 -131
rect 400 -132 401 -131
rect 401 -132 402 -131
rect 402 -132 403 -131
rect 403 -132 404 -131
rect 404 -132 405 -131
rect 405 -132 406 -131
rect 406 -132 407 -131
rect 407 -132 408 -131
rect 408 -132 409 -131
rect 409 -132 410 -131
rect 410 -132 411 -131
rect 411 -132 412 -131
rect 412 -132 413 -131
rect 413 -132 414 -131
rect 414 -132 415 -131
rect 415 -132 416 -131
rect 416 -132 417 -131
rect 417 -132 418 -131
rect 418 -132 419 -131
rect 419 -132 420 -131
rect 420 -132 421 -131
rect 421 -132 422 -131
rect 422 -132 423 -131
rect 423 -132 424 -131
rect 424 -132 425 -131
rect 425 -132 426 -131
rect 426 -132 427 -131
rect 427 -132 428 -131
rect 428 -132 429 -131
rect 429 -132 430 -131
rect 430 -132 431 -131
rect 431 -132 432 -131
rect 432 -132 433 -131
rect 433 -132 434 -131
rect 434 -132 435 -131
rect 435 -132 436 -131
rect 436 -132 437 -131
rect 437 -132 438 -131
rect 438 -132 439 -131
rect 439 -132 440 -131
rect 440 -132 441 -131
rect 441 -132 442 -131
rect 442 -132 443 -131
rect 443 -132 444 -131
rect 444 -132 445 -131
rect 445 -132 446 -131
rect 446 -132 447 -131
rect 447 -132 448 -131
rect 448 -132 449 -131
rect 449 -132 450 -131
rect 450 -132 451 -131
rect 451 -132 452 -131
rect 452 -132 453 -131
rect 453 -132 454 -131
rect 454 -132 455 -131
rect 455 -132 456 -131
rect 456 -132 457 -131
rect 457 -132 458 -131
rect 458 -132 459 -131
rect 459 -132 460 -131
rect 460 -132 461 -131
rect 461 -132 462 -131
rect 462 -132 463 -131
rect 463 -132 464 -131
rect 464 -132 465 -131
rect 465 -132 466 -131
rect 466 -132 467 -131
rect 467 -132 468 -131
rect 468 -132 469 -131
rect 469 -132 470 -131
rect 470 -132 471 -131
rect 471 -132 472 -131
rect 472 -132 473 -131
rect 473 -132 474 -131
rect 474 -132 475 -131
rect 475 -132 476 -131
rect 476 -132 477 -131
rect 477 -132 478 -131
rect 478 -132 479 -131
rect 479 -132 480 -131
rect 2 -133 3 -132
rect 3 -133 4 -132
rect 4 -133 5 -132
rect 5 -133 6 -132
rect 6 -133 7 -132
rect 7 -133 8 -132
rect 8 -133 9 -132
rect 9 -133 10 -132
rect 10 -133 11 -132
rect 11 -133 12 -132
rect 12 -133 13 -132
rect 13 -133 14 -132
rect 14 -133 15 -132
rect 15 -133 16 -132
rect 16 -133 17 -132
rect 17 -133 18 -132
rect 18 -133 19 -132
rect 19 -133 20 -132
rect 20 -133 21 -132
rect 21 -133 22 -132
rect 22 -133 23 -132
rect 23 -133 24 -132
rect 24 -133 25 -132
rect 25 -133 26 -132
rect 26 -133 27 -132
rect 27 -133 28 -132
rect 28 -133 29 -132
rect 29 -133 30 -132
rect 30 -133 31 -132
rect 31 -133 32 -132
rect 32 -133 33 -132
rect 33 -133 34 -132
rect 34 -133 35 -132
rect 35 -133 36 -132
rect 36 -133 37 -132
rect 37 -133 38 -132
rect 38 -133 39 -132
rect 39 -133 40 -132
rect 40 -133 41 -132
rect 41 -133 42 -132
rect 42 -133 43 -132
rect 43 -133 44 -132
rect 44 -133 45 -132
rect 45 -133 46 -132
rect 46 -133 47 -132
rect 47 -133 48 -132
rect 48 -133 49 -132
rect 49 -133 50 -132
rect 50 -133 51 -132
rect 51 -133 52 -132
rect 52 -133 53 -132
rect 53 -133 54 -132
rect 54 -133 55 -132
rect 55 -133 56 -132
rect 56 -133 57 -132
rect 57 -133 58 -132
rect 58 -133 59 -132
rect 59 -133 60 -132
rect 60 -133 61 -132
rect 61 -133 62 -132
rect 62 -133 63 -132
rect 63 -133 64 -132
rect 64 -133 65 -132
rect 65 -133 66 -132
rect 66 -133 67 -132
rect 67 -133 68 -132
rect 68 -133 69 -132
rect 69 -133 70 -132
rect 70 -133 71 -132
rect 71 -133 72 -132
rect 72 -133 73 -132
rect 73 -133 74 -132
rect 74 -133 75 -132
rect 75 -133 76 -132
rect 76 -133 77 -132
rect 77 -133 78 -132
rect 78 -133 79 -132
rect 79 -133 80 -132
rect 80 -133 81 -132
rect 81 -133 82 -132
rect 82 -133 83 -132
rect 83 -133 84 -132
rect 84 -133 85 -132
rect 85 -133 86 -132
rect 86 -133 87 -132
rect 87 -133 88 -132
rect 88 -133 89 -132
rect 89 -133 90 -132
rect 90 -133 91 -132
rect 91 -133 92 -132
rect 92 -133 93 -132
rect 93 -133 94 -132
rect 94 -133 95 -132
rect 95 -133 96 -132
rect 96 -133 97 -132
rect 97 -133 98 -132
rect 98 -133 99 -132
rect 99 -133 100 -132
rect 100 -133 101 -132
rect 101 -133 102 -132
rect 102 -133 103 -132
rect 103 -133 104 -132
rect 104 -133 105 -132
rect 105 -133 106 -132
rect 106 -133 107 -132
rect 107 -133 108 -132
rect 108 -133 109 -132
rect 109 -133 110 -132
rect 110 -133 111 -132
rect 111 -133 112 -132
rect 112 -133 113 -132
rect 113 -133 114 -132
rect 114 -133 115 -132
rect 115 -133 116 -132
rect 116 -133 117 -132
rect 117 -133 118 -132
rect 118 -133 119 -132
rect 119 -133 120 -132
rect 120 -133 121 -132
rect 121 -133 122 -132
rect 122 -133 123 -132
rect 123 -133 124 -132
rect 124 -133 125 -132
rect 125 -133 126 -132
rect 126 -133 127 -132
rect 127 -133 128 -132
rect 128 -133 129 -132
rect 129 -133 130 -132
rect 130 -133 131 -132
rect 131 -133 132 -132
rect 132 -133 133 -132
rect 133 -133 134 -132
rect 134 -133 135 -132
rect 135 -133 136 -132
rect 136 -133 137 -132
rect 137 -133 138 -132
rect 138 -133 139 -132
rect 139 -133 140 -132
rect 140 -133 141 -132
rect 141 -133 142 -132
rect 142 -133 143 -132
rect 143 -133 144 -132
rect 144 -133 145 -132
rect 145 -133 146 -132
rect 146 -133 147 -132
rect 147 -133 148 -132
rect 148 -133 149 -132
rect 149 -133 150 -132
rect 150 -133 151 -132
rect 151 -133 152 -132
rect 152 -133 153 -132
rect 153 -133 154 -132
rect 154 -133 155 -132
rect 155 -133 156 -132
rect 156 -133 157 -132
rect 157 -133 158 -132
rect 158 -133 159 -132
rect 159 -133 160 -132
rect 160 -133 161 -132
rect 161 -133 162 -132
rect 162 -133 163 -132
rect 163 -133 164 -132
rect 164 -133 165 -132
rect 165 -133 166 -132
rect 166 -133 167 -132
rect 167 -133 168 -132
rect 168 -133 169 -132
rect 169 -133 170 -132
rect 170 -133 171 -132
rect 171 -133 172 -132
rect 172 -133 173 -132
rect 173 -133 174 -132
rect 174 -133 175 -132
rect 175 -133 176 -132
rect 176 -133 177 -132
rect 177 -133 178 -132
rect 178 -133 179 -132
rect 179 -133 180 -132
rect 180 -133 181 -132
rect 181 -133 182 -132
rect 182 -133 183 -132
rect 183 -133 184 -132
rect 184 -133 185 -132
rect 185 -133 186 -132
rect 186 -133 187 -132
rect 187 -133 188 -132
rect 188 -133 189 -132
rect 189 -133 190 -132
rect 190 -133 191 -132
rect 191 -133 192 -132
rect 192 -133 193 -132
rect 193 -133 194 -132
rect 194 -133 195 -132
rect 195 -133 196 -132
rect 196 -133 197 -132
rect 197 -133 198 -132
rect 198 -133 199 -132
rect 199 -133 200 -132
rect 200 -133 201 -132
rect 201 -133 202 -132
rect 202 -133 203 -132
rect 203 -133 204 -132
rect 204 -133 205 -132
rect 205 -133 206 -132
rect 206 -133 207 -132
rect 207 -133 208 -132
rect 208 -133 209 -132
rect 209 -133 210 -132
rect 210 -133 211 -132
rect 211 -133 212 -132
rect 212 -133 213 -132
rect 213 -133 214 -132
rect 214 -133 215 -132
rect 215 -133 216 -132
rect 216 -133 217 -132
rect 217 -133 218 -132
rect 218 -133 219 -132
rect 219 -133 220 -132
rect 220 -133 221 -132
rect 221 -133 222 -132
rect 222 -133 223 -132
rect 223 -133 224 -132
rect 224 -133 225 -132
rect 225 -133 226 -132
rect 226 -133 227 -132
rect 227 -133 228 -132
rect 228 -133 229 -132
rect 229 -133 230 -132
rect 230 -133 231 -132
rect 231 -133 232 -132
rect 232 -133 233 -132
rect 233 -133 234 -132
rect 234 -133 235 -132
rect 235 -133 236 -132
rect 236 -133 237 -132
rect 237 -133 238 -132
rect 238 -133 239 -132
rect 239 -133 240 -132
rect 240 -133 241 -132
rect 241 -133 242 -132
rect 242 -133 243 -132
rect 243 -133 244 -132
rect 244 -133 245 -132
rect 245 -133 246 -132
rect 246 -133 247 -132
rect 247 -133 248 -132
rect 248 -133 249 -132
rect 249 -133 250 -132
rect 250 -133 251 -132
rect 251 -133 252 -132
rect 252 -133 253 -132
rect 253 -133 254 -132
rect 254 -133 255 -132
rect 255 -133 256 -132
rect 256 -133 257 -132
rect 257 -133 258 -132
rect 258 -133 259 -132
rect 259 -133 260 -132
rect 260 -133 261 -132
rect 261 -133 262 -132
rect 262 -133 263 -132
rect 263 -133 264 -132
rect 264 -133 265 -132
rect 265 -133 266 -132
rect 266 -133 267 -132
rect 267 -133 268 -132
rect 268 -133 269 -132
rect 269 -133 270 -132
rect 270 -133 271 -132
rect 271 -133 272 -132
rect 272 -133 273 -132
rect 273 -133 274 -132
rect 274 -133 275 -132
rect 275 -133 276 -132
rect 276 -133 277 -132
rect 277 -133 278 -132
rect 278 -133 279 -132
rect 279 -133 280 -132
rect 280 -133 281 -132
rect 281 -133 282 -132
rect 282 -133 283 -132
rect 283 -133 284 -132
rect 284 -133 285 -132
rect 285 -133 286 -132
rect 286 -133 287 -132
rect 287 -133 288 -132
rect 288 -133 289 -132
rect 289 -133 290 -132
rect 290 -133 291 -132
rect 291 -133 292 -132
rect 292 -133 293 -132
rect 293 -133 294 -132
rect 294 -133 295 -132
rect 295 -133 296 -132
rect 296 -133 297 -132
rect 297 -133 298 -132
rect 298 -133 299 -132
rect 299 -133 300 -132
rect 300 -133 301 -132
rect 301 -133 302 -132
rect 302 -133 303 -132
rect 303 -133 304 -132
rect 304 -133 305 -132
rect 305 -133 306 -132
rect 306 -133 307 -132
rect 307 -133 308 -132
rect 308 -133 309 -132
rect 309 -133 310 -132
rect 310 -133 311 -132
rect 311 -133 312 -132
rect 312 -133 313 -132
rect 313 -133 314 -132
rect 314 -133 315 -132
rect 315 -133 316 -132
rect 316 -133 317 -132
rect 317 -133 318 -132
rect 318 -133 319 -132
rect 319 -133 320 -132
rect 320 -133 321 -132
rect 321 -133 322 -132
rect 322 -133 323 -132
rect 323 -133 324 -132
rect 324 -133 325 -132
rect 325 -133 326 -132
rect 326 -133 327 -132
rect 327 -133 328 -132
rect 328 -133 329 -132
rect 329 -133 330 -132
rect 330 -133 331 -132
rect 331 -133 332 -132
rect 332 -133 333 -132
rect 333 -133 334 -132
rect 334 -133 335 -132
rect 335 -133 336 -132
rect 336 -133 337 -132
rect 337 -133 338 -132
rect 338 -133 339 -132
rect 339 -133 340 -132
rect 340 -133 341 -132
rect 341 -133 342 -132
rect 342 -133 343 -132
rect 343 -133 344 -132
rect 344 -133 345 -132
rect 345 -133 346 -132
rect 346 -133 347 -132
rect 347 -133 348 -132
rect 348 -133 349 -132
rect 349 -133 350 -132
rect 350 -133 351 -132
rect 351 -133 352 -132
rect 352 -133 353 -132
rect 353 -133 354 -132
rect 354 -133 355 -132
rect 355 -133 356 -132
rect 356 -133 357 -132
rect 357 -133 358 -132
rect 358 -133 359 -132
rect 359 -133 360 -132
rect 360 -133 361 -132
rect 361 -133 362 -132
rect 362 -133 363 -132
rect 363 -133 364 -132
rect 364 -133 365 -132
rect 365 -133 366 -132
rect 366 -133 367 -132
rect 367 -133 368 -132
rect 368 -133 369 -132
rect 369 -133 370 -132
rect 370 -133 371 -132
rect 371 -133 372 -132
rect 372 -133 373 -132
rect 373 -133 374 -132
rect 374 -133 375 -132
rect 375 -133 376 -132
rect 376 -133 377 -132
rect 377 -133 378 -132
rect 378 -133 379 -132
rect 379 -133 380 -132
rect 380 -133 381 -132
rect 381 -133 382 -132
rect 382 -133 383 -132
rect 383 -133 384 -132
rect 384 -133 385 -132
rect 385 -133 386 -132
rect 386 -133 387 -132
rect 387 -133 388 -132
rect 388 -133 389 -132
rect 389 -133 390 -132
rect 390 -133 391 -132
rect 391 -133 392 -132
rect 392 -133 393 -132
rect 393 -133 394 -132
rect 394 -133 395 -132
rect 395 -133 396 -132
rect 396 -133 397 -132
rect 397 -133 398 -132
rect 398 -133 399 -132
rect 399 -133 400 -132
rect 400 -133 401 -132
rect 401 -133 402 -132
rect 402 -133 403 -132
rect 403 -133 404 -132
rect 404 -133 405 -132
rect 405 -133 406 -132
rect 406 -133 407 -132
rect 407 -133 408 -132
rect 408 -133 409 -132
rect 409 -133 410 -132
rect 410 -133 411 -132
rect 411 -133 412 -132
rect 412 -133 413 -132
rect 413 -133 414 -132
rect 414 -133 415 -132
rect 415 -133 416 -132
rect 416 -133 417 -132
rect 417 -133 418 -132
rect 418 -133 419 -132
rect 419 -133 420 -132
rect 420 -133 421 -132
rect 421 -133 422 -132
rect 422 -133 423 -132
rect 423 -133 424 -132
rect 424 -133 425 -132
rect 425 -133 426 -132
rect 426 -133 427 -132
rect 427 -133 428 -132
rect 428 -133 429 -132
rect 429 -133 430 -132
rect 430 -133 431 -132
rect 431 -133 432 -132
rect 432 -133 433 -132
rect 433 -133 434 -132
rect 434 -133 435 -132
rect 435 -133 436 -132
rect 436 -133 437 -132
rect 437 -133 438 -132
rect 438 -133 439 -132
rect 439 -133 440 -132
rect 440 -133 441 -132
rect 441 -133 442 -132
rect 442 -133 443 -132
rect 443 -133 444 -132
rect 444 -133 445 -132
rect 445 -133 446 -132
rect 446 -133 447 -132
rect 447 -133 448 -132
rect 448 -133 449 -132
rect 449 -133 450 -132
rect 450 -133 451 -132
rect 451 -133 452 -132
rect 452 -133 453 -132
rect 453 -133 454 -132
rect 454 -133 455 -132
rect 455 -133 456 -132
rect 456 -133 457 -132
rect 457 -133 458 -132
rect 458 -133 459 -132
rect 459 -133 460 -132
rect 460 -133 461 -132
rect 461 -133 462 -132
rect 462 -133 463 -132
rect 463 -133 464 -132
rect 464 -133 465 -132
rect 465 -133 466 -132
rect 466 -133 467 -132
rect 467 -133 468 -132
rect 468 -133 469 -132
rect 469 -133 470 -132
rect 470 -133 471 -132
rect 471 -133 472 -132
rect 472 -133 473 -132
rect 473 -133 474 -132
rect 474 -133 475 -132
rect 475 -133 476 -132
rect 476 -133 477 -132
rect 477 -133 478 -132
rect 478 -133 479 -132
rect 479 -133 480 -132
rect 2 -134 3 -133
rect 3 -134 4 -133
rect 4 -134 5 -133
rect 5 -134 6 -133
rect 6 -134 7 -133
rect 7 -134 8 -133
rect 8 -134 9 -133
rect 9 -134 10 -133
rect 10 -134 11 -133
rect 11 -134 12 -133
rect 12 -134 13 -133
rect 13 -134 14 -133
rect 14 -134 15 -133
rect 15 -134 16 -133
rect 16 -134 17 -133
rect 17 -134 18 -133
rect 18 -134 19 -133
rect 19 -134 20 -133
rect 20 -134 21 -133
rect 21 -134 22 -133
rect 22 -134 23 -133
rect 23 -134 24 -133
rect 24 -134 25 -133
rect 25 -134 26 -133
rect 26 -134 27 -133
rect 27 -134 28 -133
rect 28 -134 29 -133
rect 29 -134 30 -133
rect 30 -134 31 -133
rect 31 -134 32 -133
rect 32 -134 33 -133
rect 33 -134 34 -133
rect 34 -134 35 -133
rect 35 -134 36 -133
rect 36 -134 37 -133
rect 37 -134 38 -133
rect 38 -134 39 -133
rect 39 -134 40 -133
rect 40 -134 41 -133
rect 41 -134 42 -133
rect 42 -134 43 -133
rect 43 -134 44 -133
rect 44 -134 45 -133
rect 45 -134 46 -133
rect 46 -134 47 -133
rect 47 -134 48 -133
rect 48 -134 49 -133
rect 49 -134 50 -133
rect 50 -134 51 -133
rect 51 -134 52 -133
rect 52 -134 53 -133
rect 53 -134 54 -133
rect 54 -134 55 -133
rect 55 -134 56 -133
rect 56 -134 57 -133
rect 57 -134 58 -133
rect 58 -134 59 -133
rect 59 -134 60 -133
rect 60 -134 61 -133
rect 61 -134 62 -133
rect 62 -134 63 -133
rect 63 -134 64 -133
rect 64 -134 65 -133
rect 65 -134 66 -133
rect 66 -134 67 -133
rect 67 -134 68 -133
rect 68 -134 69 -133
rect 69 -134 70 -133
rect 70 -134 71 -133
rect 71 -134 72 -133
rect 72 -134 73 -133
rect 73 -134 74 -133
rect 74 -134 75 -133
rect 75 -134 76 -133
rect 76 -134 77 -133
rect 77 -134 78 -133
rect 78 -134 79 -133
rect 79 -134 80 -133
rect 80 -134 81 -133
rect 81 -134 82 -133
rect 82 -134 83 -133
rect 83 -134 84 -133
rect 84 -134 85 -133
rect 85 -134 86 -133
rect 86 -134 87 -133
rect 87 -134 88 -133
rect 88 -134 89 -133
rect 89 -134 90 -133
rect 90 -134 91 -133
rect 91 -134 92 -133
rect 92 -134 93 -133
rect 93 -134 94 -133
rect 94 -134 95 -133
rect 95 -134 96 -133
rect 96 -134 97 -133
rect 97 -134 98 -133
rect 98 -134 99 -133
rect 99 -134 100 -133
rect 100 -134 101 -133
rect 101 -134 102 -133
rect 102 -134 103 -133
rect 103 -134 104 -133
rect 104 -134 105 -133
rect 105 -134 106 -133
rect 106 -134 107 -133
rect 107 -134 108 -133
rect 108 -134 109 -133
rect 109 -134 110 -133
rect 110 -134 111 -133
rect 111 -134 112 -133
rect 112 -134 113 -133
rect 113 -134 114 -133
rect 114 -134 115 -133
rect 115 -134 116 -133
rect 116 -134 117 -133
rect 117 -134 118 -133
rect 118 -134 119 -133
rect 119 -134 120 -133
rect 120 -134 121 -133
rect 121 -134 122 -133
rect 122 -134 123 -133
rect 123 -134 124 -133
rect 124 -134 125 -133
rect 125 -134 126 -133
rect 126 -134 127 -133
rect 127 -134 128 -133
rect 128 -134 129 -133
rect 129 -134 130 -133
rect 130 -134 131 -133
rect 131 -134 132 -133
rect 132 -134 133 -133
rect 133 -134 134 -133
rect 134 -134 135 -133
rect 135 -134 136 -133
rect 136 -134 137 -133
rect 137 -134 138 -133
rect 138 -134 139 -133
rect 139 -134 140 -133
rect 140 -134 141 -133
rect 141 -134 142 -133
rect 142 -134 143 -133
rect 143 -134 144 -133
rect 144 -134 145 -133
rect 145 -134 146 -133
rect 146 -134 147 -133
rect 147 -134 148 -133
rect 148 -134 149 -133
rect 149 -134 150 -133
rect 150 -134 151 -133
rect 151 -134 152 -133
rect 152 -134 153 -133
rect 153 -134 154 -133
rect 154 -134 155 -133
rect 155 -134 156 -133
rect 156 -134 157 -133
rect 157 -134 158 -133
rect 158 -134 159 -133
rect 159 -134 160 -133
rect 160 -134 161 -133
rect 161 -134 162 -133
rect 162 -134 163 -133
rect 163 -134 164 -133
rect 164 -134 165 -133
rect 165 -134 166 -133
rect 166 -134 167 -133
rect 167 -134 168 -133
rect 168 -134 169 -133
rect 169 -134 170 -133
rect 170 -134 171 -133
rect 171 -134 172 -133
rect 172 -134 173 -133
rect 173 -134 174 -133
rect 174 -134 175 -133
rect 175 -134 176 -133
rect 176 -134 177 -133
rect 177 -134 178 -133
rect 178 -134 179 -133
rect 179 -134 180 -133
rect 180 -134 181 -133
rect 181 -134 182 -133
rect 182 -134 183 -133
rect 183 -134 184 -133
rect 184 -134 185 -133
rect 185 -134 186 -133
rect 186 -134 187 -133
rect 187 -134 188 -133
rect 188 -134 189 -133
rect 189 -134 190 -133
rect 190 -134 191 -133
rect 191 -134 192 -133
rect 192 -134 193 -133
rect 193 -134 194 -133
rect 194 -134 195 -133
rect 195 -134 196 -133
rect 196 -134 197 -133
rect 197 -134 198 -133
rect 198 -134 199 -133
rect 199 -134 200 -133
rect 200 -134 201 -133
rect 201 -134 202 -133
rect 202 -134 203 -133
rect 203 -134 204 -133
rect 204 -134 205 -133
rect 205 -134 206 -133
rect 206 -134 207 -133
rect 207 -134 208 -133
rect 208 -134 209 -133
rect 209 -134 210 -133
rect 210 -134 211 -133
rect 211 -134 212 -133
rect 212 -134 213 -133
rect 213 -134 214 -133
rect 214 -134 215 -133
rect 215 -134 216 -133
rect 216 -134 217 -133
rect 217 -134 218 -133
rect 218 -134 219 -133
rect 219 -134 220 -133
rect 220 -134 221 -133
rect 221 -134 222 -133
rect 222 -134 223 -133
rect 223 -134 224 -133
rect 224 -134 225 -133
rect 225 -134 226 -133
rect 226 -134 227 -133
rect 227 -134 228 -133
rect 228 -134 229 -133
rect 229 -134 230 -133
rect 230 -134 231 -133
rect 231 -134 232 -133
rect 232 -134 233 -133
rect 233 -134 234 -133
rect 234 -134 235 -133
rect 235 -134 236 -133
rect 236 -134 237 -133
rect 237 -134 238 -133
rect 238 -134 239 -133
rect 239 -134 240 -133
rect 240 -134 241 -133
rect 241 -134 242 -133
rect 242 -134 243 -133
rect 243 -134 244 -133
rect 244 -134 245 -133
rect 245 -134 246 -133
rect 246 -134 247 -133
rect 247 -134 248 -133
rect 248 -134 249 -133
rect 249 -134 250 -133
rect 250 -134 251 -133
rect 251 -134 252 -133
rect 252 -134 253 -133
rect 253 -134 254 -133
rect 254 -134 255 -133
rect 255 -134 256 -133
rect 256 -134 257 -133
rect 257 -134 258 -133
rect 258 -134 259 -133
rect 259 -134 260 -133
rect 260 -134 261 -133
rect 261 -134 262 -133
rect 262 -134 263 -133
rect 263 -134 264 -133
rect 264 -134 265 -133
rect 265 -134 266 -133
rect 266 -134 267 -133
rect 267 -134 268 -133
rect 268 -134 269 -133
rect 269 -134 270 -133
rect 270 -134 271 -133
rect 271 -134 272 -133
rect 272 -134 273 -133
rect 273 -134 274 -133
rect 274 -134 275 -133
rect 275 -134 276 -133
rect 276 -134 277 -133
rect 277 -134 278 -133
rect 278 -134 279 -133
rect 279 -134 280 -133
rect 280 -134 281 -133
rect 281 -134 282 -133
rect 282 -134 283 -133
rect 283 -134 284 -133
rect 284 -134 285 -133
rect 285 -134 286 -133
rect 286 -134 287 -133
rect 287 -134 288 -133
rect 288 -134 289 -133
rect 289 -134 290 -133
rect 290 -134 291 -133
rect 291 -134 292 -133
rect 292 -134 293 -133
rect 293 -134 294 -133
rect 294 -134 295 -133
rect 295 -134 296 -133
rect 296 -134 297 -133
rect 297 -134 298 -133
rect 298 -134 299 -133
rect 299 -134 300 -133
rect 300 -134 301 -133
rect 301 -134 302 -133
rect 302 -134 303 -133
rect 303 -134 304 -133
rect 304 -134 305 -133
rect 305 -134 306 -133
rect 306 -134 307 -133
rect 307 -134 308 -133
rect 308 -134 309 -133
rect 309 -134 310 -133
rect 310 -134 311 -133
rect 311 -134 312 -133
rect 312 -134 313 -133
rect 313 -134 314 -133
rect 314 -134 315 -133
rect 315 -134 316 -133
rect 316 -134 317 -133
rect 317 -134 318 -133
rect 318 -134 319 -133
rect 319 -134 320 -133
rect 320 -134 321 -133
rect 321 -134 322 -133
rect 322 -134 323 -133
rect 323 -134 324 -133
rect 324 -134 325 -133
rect 325 -134 326 -133
rect 326 -134 327 -133
rect 327 -134 328 -133
rect 328 -134 329 -133
rect 329 -134 330 -133
rect 330 -134 331 -133
rect 331 -134 332 -133
rect 332 -134 333 -133
rect 333 -134 334 -133
rect 334 -134 335 -133
rect 335 -134 336 -133
rect 336 -134 337 -133
rect 337 -134 338 -133
rect 338 -134 339 -133
rect 339 -134 340 -133
rect 340 -134 341 -133
rect 341 -134 342 -133
rect 342 -134 343 -133
rect 343 -134 344 -133
rect 344 -134 345 -133
rect 345 -134 346 -133
rect 346 -134 347 -133
rect 347 -134 348 -133
rect 348 -134 349 -133
rect 349 -134 350 -133
rect 350 -134 351 -133
rect 351 -134 352 -133
rect 352 -134 353 -133
rect 353 -134 354 -133
rect 354 -134 355 -133
rect 355 -134 356 -133
rect 356 -134 357 -133
rect 357 -134 358 -133
rect 358 -134 359 -133
rect 359 -134 360 -133
rect 360 -134 361 -133
rect 361 -134 362 -133
rect 362 -134 363 -133
rect 363 -134 364 -133
rect 364 -134 365 -133
rect 365 -134 366 -133
rect 366 -134 367 -133
rect 367 -134 368 -133
rect 368 -134 369 -133
rect 369 -134 370 -133
rect 370 -134 371 -133
rect 371 -134 372 -133
rect 372 -134 373 -133
rect 373 -134 374 -133
rect 374 -134 375 -133
rect 375 -134 376 -133
rect 376 -134 377 -133
rect 377 -134 378 -133
rect 378 -134 379 -133
rect 379 -134 380 -133
rect 380 -134 381 -133
rect 381 -134 382 -133
rect 382 -134 383 -133
rect 383 -134 384 -133
rect 384 -134 385 -133
rect 385 -134 386 -133
rect 386 -134 387 -133
rect 387 -134 388 -133
rect 388 -134 389 -133
rect 389 -134 390 -133
rect 390 -134 391 -133
rect 391 -134 392 -133
rect 392 -134 393 -133
rect 393 -134 394 -133
rect 394 -134 395 -133
rect 395 -134 396 -133
rect 396 -134 397 -133
rect 397 -134 398 -133
rect 398 -134 399 -133
rect 399 -134 400 -133
rect 400 -134 401 -133
rect 401 -134 402 -133
rect 402 -134 403 -133
rect 403 -134 404 -133
rect 404 -134 405 -133
rect 405 -134 406 -133
rect 406 -134 407 -133
rect 407 -134 408 -133
rect 408 -134 409 -133
rect 409 -134 410 -133
rect 410 -134 411 -133
rect 411 -134 412 -133
rect 412 -134 413 -133
rect 413 -134 414 -133
rect 414 -134 415 -133
rect 415 -134 416 -133
rect 416 -134 417 -133
rect 417 -134 418 -133
rect 418 -134 419 -133
rect 419 -134 420 -133
rect 420 -134 421 -133
rect 421 -134 422 -133
rect 422 -134 423 -133
rect 423 -134 424 -133
rect 424 -134 425 -133
rect 425 -134 426 -133
rect 426 -134 427 -133
rect 427 -134 428 -133
rect 428 -134 429 -133
rect 429 -134 430 -133
rect 430 -134 431 -133
rect 431 -134 432 -133
rect 432 -134 433 -133
rect 433 -134 434 -133
rect 434 -134 435 -133
rect 435 -134 436 -133
rect 436 -134 437 -133
rect 437 -134 438 -133
rect 438 -134 439 -133
rect 439 -134 440 -133
rect 440 -134 441 -133
rect 441 -134 442 -133
rect 442 -134 443 -133
rect 443 -134 444 -133
rect 444 -134 445 -133
rect 445 -134 446 -133
rect 446 -134 447 -133
rect 447 -134 448 -133
rect 448 -134 449 -133
rect 449 -134 450 -133
rect 450 -134 451 -133
rect 451 -134 452 -133
rect 452 -134 453 -133
rect 453 -134 454 -133
rect 454 -134 455 -133
rect 455 -134 456 -133
rect 456 -134 457 -133
rect 457 -134 458 -133
rect 458 -134 459 -133
rect 459 -134 460 -133
rect 460 -134 461 -133
rect 461 -134 462 -133
rect 462 -134 463 -133
rect 463 -134 464 -133
rect 464 -134 465 -133
rect 465 -134 466 -133
rect 466 -134 467 -133
rect 467 -134 468 -133
rect 468 -134 469 -133
rect 469 -134 470 -133
rect 470 -134 471 -133
rect 471 -134 472 -133
rect 472 -134 473 -133
rect 473 -134 474 -133
rect 474 -134 475 -133
rect 475 -134 476 -133
rect 476 -134 477 -133
rect 477 -134 478 -133
rect 478 -134 479 -133
rect 479 -134 480 -133
rect 2 -157 3 -156
rect 3 -157 4 -156
rect 4 -157 5 -156
rect 5 -157 6 -156
rect 6 -157 7 -156
rect 7 -157 8 -156
rect 8 -157 9 -156
rect 9 -157 10 -156
rect 10 -157 11 -156
rect 11 -157 12 -156
rect 12 -157 13 -156
rect 13 -157 14 -156
rect 14 -157 15 -156
rect 15 -157 16 -156
rect 16 -157 17 -156
rect 17 -157 18 -156
rect 18 -157 19 -156
rect 19 -157 20 -156
rect 20 -157 21 -156
rect 21 -157 22 -156
rect 22 -157 23 -156
rect 23 -157 24 -156
rect 24 -157 25 -156
rect 25 -157 26 -156
rect 26 -157 27 -156
rect 27 -157 28 -156
rect 28 -157 29 -156
rect 29 -157 30 -156
rect 30 -157 31 -156
rect 31 -157 32 -156
rect 32 -157 33 -156
rect 33 -157 34 -156
rect 34 -157 35 -156
rect 35 -157 36 -156
rect 36 -157 37 -156
rect 37 -157 38 -156
rect 38 -157 39 -156
rect 39 -157 40 -156
rect 40 -157 41 -156
rect 41 -157 42 -156
rect 42 -157 43 -156
rect 43 -157 44 -156
rect 44 -157 45 -156
rect 45 -157 46 -156
rect 46 -157 47 -156
rect 47 -157 48 -156
rect 48 -157 49 -156
rect 49 -157 50 -156
rect 50 -157 51 -156
rect 51 -157 52 -156
rect 52 -157 53 -156
rect 53 -157 54 -156
rect 54 -157 55 -156
rect 55 -157 56 -156
rect 56 -157 57 -156
rect 57 -157 58 -156
rect 58 -157 59 -156
rect 59 -157 60 -156
rect 60 -157 61 -156
rect 61 -157 62 -156
rect 62 -157 63 -156
rect 63 -157 64 -156
rect 64 -157 65 -156
rect 65 -157 66 -156
rect 66 -157 67 -156
rect 67 -157 68 -156
rect 68 -157 69 -156
rect 69 -157 70 -156
rect 70 -157 71 -156
rect 71 -157 72 -156
rect 72 -157 73 -156
rect 73 -157 74 -156
rect 74 -157 75 -156
rect 75 -157 76 -156
rect 76 -157 77 -156
rect 77 -157 78 -156
rect 78 -157 79 -156
rect 79 -157 80 -156
rect 80 -157 81 -156
rect 81 -157 82 -156
rect 82 -157 83 -156
rect 83 -157 84 -156
rect 84 -157 85 -156
rect 85 -157 86 -156
rect 86 -157 87 -156
rect 87 -157 88 -156
rect 88 -157 89 -156
rect 89 -157 90 -156
rect 90 -157 91 -156
rect 91 -157 92 -156
rect 92 -157 93 -156
rect 93 -157 94 -156
rect 94 -157 95 -156
rect 95 -157 96 -156
rect 96 -157 97 -156
rect 97 -157 98 -156
rect 98 -157 99 -156
rect 99 -157 100 -156
rect 100 -157 101 -156
rect 101 -157 102 -156
rect 102 -157 103 -156
rect 103 -157 104 -156
rect 104 -157 105 -156
rect 105 -157 106 -156
rect 106 -157 107 -156
rect 107 -157 108 -156
rect 108 -157 109 -156
rect 109 -157 110 -156
rect 110 -157 111 -156
rect 111 -157 112 -156
rect 112 -157 113 -156
rect 113 -157 114 -156
rect 114 -157 115 -156
rect 115 -157 116 -156
rect 116 -157 117 -156
rect 117 -157 118 -156
rect 118 -157 119 -156
rect 119 -157 120 -156
rect 120 -157 121 -156
rect 121 -157 122 -156
rect 122 -157 123 -156
rect 123 -157 124 -156
rect 124 -157 125 -156
rect 125 -157 126 -156
rect 126 -157 127 -156
rect 127 -157 128 -156
rect 128 -157 129 -156
rect 129 -157 130 -156
rect 130 -157 131 -156
rect 131 -157 132 -156
rect 132 -157 133 -156
rect 133 -157 134 -156
rect 134 -157 135 -156
rect 135 -157 136 -156
rect 136 -157 137 -156
rect 137 -157 138 -156
rect 138 -157 139 -156
rect 139 -157 140 -156
rect 140 -157 141 -156
rect 141 -157 142 -156
rect 142 -157 143 -156
rect 143 -157 144 -156
rect 144 -157 145 -156
rect 145 -157 146 -156
rect 146 -157 147 -156
rect 147 -157 148 -156
rect 148 -157 149 -156
rect 149 -157 150 -156
rect 150 -157 151 -156
rect 151 -157 152 -156
rect 152 -157 153 -156
rect 153 -157 154 -156
rect 154 -157 155 -156
rect 155 -157 156 -156
rect 156 -157 157 -156
rect 157 -157 158 -156
rect 158 -157 159 -156
rect 159 -157 160 -156
rect 160 -157 161 -156
rect 161 -157 162 -156
rect 162 -157 163 -156
rect 163 -157 164 -156
rect 164 -157 165 -156
rect 165 -157 166 -156
rect 166 -157 167 -156
rect 167 -157 168 -156
rect 168 -157 169 -156
rect 169 -157 170 -156
rect 170 -157 171 -156
rect 171 -157 172 -156
rect 172 -157 173 -156
rect 173 -157 174 -156
rect 174 -157 175 -156
rect 175 -157 176 -156
rect 176 -157 177 -156
rect 177 -157 178 -156
rect 178 -157 179 -156
rect 179 -157 180 -156
rect 180 -157 181 -156
rect 181 -157 182 -156
rect 182 -157 183 -156
rect 183 -157 184 -156
rect 184 -157 185 -156
rect 185 -157 186 -156
rect 186 -157 187 -156
rect 187 -157 188 -156
rect 188 -157 189 -156
rect 189 -157 190 -156
rect 190 -157 191 -156
rect 191 -157 192 -156
rect 192 -157 193 -156
rect 193 -157 194 -156
rect 194 -157 195 -156
rect 195 -157 196 -156
rect 196 -157 197 -156
rect 197 -157 198 -156
rect 198 -157 199 -156
rect 199 -157 200 -156
rect 200 -157 201 -156
rect 201 -157 202 -156
rect 202 -157 203 -156
rect 203 -157 204 -156
rect 204 -157 205 -156
rect 205 -157 206 -156
rect 206 -157 207 -156
rect 207 -157 208 -156
rect 208 -157 209 -156
rect 209 -157 210 -156
rect 210 -157 211 -156
rect 211 -157 212 -156
rect 212 -157 213 -156
rect 213 -157 214 -156
rect 214 -157 215 -156
rect 215 -157 216 -156
rect 216 -157 217 -156
rect 217 -157 218 -156
rect 218 -157 219 -156
rect 219 -157 220 -156
rect 220 -157 221 -156
rect 221 -157 222 -156
rect 222 -157 223 -156
rect 223 -157 224 -156
rect 224 -157 225 -156
rect 225 -157 226 -156
rect 226 -157 227 -156
rect 227 -157 228 -156
rect 228 -157 229 -156
rect 229 -157 230 -156
rect 230 -157 231 -156
rect 231 -157 232 -156
rect 232 -157 233 -156
rect 233 -157 234 -156
rect 234 -157 235 -156
rect 235 -157 236 -156
rect 236 -157 237 -156
rect 237 -157 238 -156
rect 238 -157 239 -156
rect 239 -157 240 -156
rect 240 -157 241 -156
rect 241 -157 242 -156
rect 242 -157 243 -156
rect 243 -157 244 -156
rect 244 -157 245 -156
rect 245 -157 246 -156
rect 246 -157 247 -156
rect 247 -157 248 -156
rect 248 -157 249 -156
rect 249 -157 250 -156
rect 250 -157 251 -156
rect 251 -157 252 -156
rect 252 -157 253 -156
rect 253 -157 254 -156
rect 254 -157 255 -156
rect 255 -157 256 -156
rect 256 -157 257 -156
rect 257 -157 258 -156
rect 258 -157 259 -156
rect 259 -157 260 -156
rect 260 -157 261 -156
rect 261 -157 262 -156
rect 262 -157 263 -156
rect 263 -157 264 -156
rect 264 -157 265 -156
rect 265 -157 266 -156
rect 266 -157 267 -156
rect 267 -157 268 -156
rect 268 -157 269 -156
rect 269 -157 270 -156
rect 270 -157 271 -156
rect 271 -157 272 -156
rect 272 -157 273 -156
rect 273 -157 274 -156
rect 274 -157 275 -156
rect 275 -157 276 -156
rect 276 -157 277 -156
rect 277 -157 278 -156
rect 278 -157 279 -156
rect 279 -157 280 -156
rect 280 -157 281 -156
rect 281 -157 282 -156
rect 282 -157 283 -156
rect 283 -157 284 -156
rect 284 -157 285 -156
rect 285 -157 286 -156
rect 286 -157 287 -156
rect 287 -157 288 -156
rect 288 -157 289 -156
rect 289 -157 290 -156
rect 290 -157 291 -156
rect 291 -157 292 -156
rect 292 -157 293 -156
rect 293 -157 294 -156
rect 294 -157 295 -156
rect 295 -157 296 -156
rect 296 -157 297 -156
rect 297 -157 298 -156
rect 298 -157 299 -156
rect 299 -157 300 -156
rect 300 -157 301 -156
rect 301 -157 302 -156
rect 302 -157 303 -156
rect 303 -157 304 -156
rect 304 -157 305 -156
rect 305 -157 306 -156
rect 306 -157 307 -156
rect 307 -157 308 -156
rect 308 -157 309 -156
rect 309 -157 310 -156
rect 310 -157 311 -156
rect 311 -157 312 -156
rect 312 -157 313 -156
rect 313 -157 314 -156
rect 314 -157 315 -156
rect 315 -157 316 -156
rect 316 -157 317 -156
rect 317 -157 318 -156
rect 318 -157 319 -156
rect 319 -157 320 -156
rect 320 -157 321 -156
rect 321 -157 322 -156
rect 322 -157 323 -156
rect 323 -157 324 -156
rect 324 -157 325 -156
rect 325 -157 326 -156
rect 326 -157 327 -156
rect 327 -157 328 -156
rect 328 -157 329 -156
rect 329 -157 330 -156
rect 330 -157 331 -156
rect 331 -157 332 -156
rect 332 -157 333 -156
rect 333 -157 334 -156
rect 334 -157 335 -156
rect 335 -157 336 -156
rect 336 -157 337 -156
rect 337 -157 338 -156
rect 338 -157 339 -156
rect 339 -157 340 -156
rect 340 -157 341 -156
rect 341 -157 342 -156
rect 342 -157 343 -156
rect 343 -157 344 -156
rect 344 -157 345 -156
rect 345 -157 346 -156
rect 346 -157 347 -156
rect 347 -157 348 -156
rect 348 -157 349 -156
rect 349 -157 350 -156
rect 350 -157 351 -156
rect 351 -157 352 -156
rect 352 -157 353 -156
rect 353 -157 354 -156
rect 354 -157 355 -156
rect 355 -157 356 -156
rect 356 -157 357 -156
rect 357 -157 358 -156
rect 358 -157 359 -156
rect 359 -157 360 -156
rect 360 -157 361 -156
rect 361 -157 362 -156
rect 362 -157 363 -156
rect 363 -157 364 -156
rect 364 -157 365 -156
rect 365 -157 366 -156
rect 366 -157 367 -156
rect 367 -157 368 -156
rect 368 -157 369 -156
rect 369 -157 370 -156
rect 370 -157 371 -156
rect 371 -157 372 -156
rect 372 -157 373 -156
rect 373 -157 374 -156
rect 374 -157 375 -156
rect 375 -157 376 -156
rect 376 -157 377 -156
rect 377 -157 378 -156
rect 378 -157 379 -156
rect 379 -157 380 -156
rect 380 -157 381 -156
rect 381 -157 382 -156
rect 382 -157 383 -156
rect 383 -157 384 -156
rect 384 -157 385 -156
rect 385 -157 386 -156
rect 386 -157 387 -156
rect 387 -157 388 -156
rect 388 -157 389 -156
rect 389 -157 390 -156
rect 390 -157 391 -156
rect 391 -157 392 -156
rect 392 -157 393 -156
rect 393 -157 394 -156
rect 394 -157 395 -156
rect 395 -157 396 -156
rect 396 -157 397 -156
rect 397 -157 398 -156
rect 398 -157 399 -156
rect 399 -157 400 -156
rect 400 -157 401 -156
rect 401 -157 402 -156
rect 402 -157 403 -156
rect 403 -157 404 -156
rect 404 -157 405 -156
rect 405 -157 406 -156
rect 406 -157 407 -156
rect 407 -157 408 -156
rect 408 -157 409 -156
rect 409 -157 410 -156
rect 410 -157 411 -156
rect 411 -157 412 -156
rect 412 -157 413 -156
rect 413 -157 414 -156
rect 414 -157 415 -156
rect 415 -157 416 -156
rect 416 -157 417 -156
rect 417 -157 418 -156
rect 418 -157 419 -156
rect 419 -157 420 -156
rect 420 -157 421 -156
rect 421 -157 422 -156
rect 422 -157 423 -156
rect 423 -157 424 -156
rect 424 -157 425 -156
rect 425 -157 426 -156
rect 426 -157 427 -156
rect 427 -157 428 -156
rect 428 -157 429 -156
rect 429 -157 430 -156
rect 430 -157 431 -156
rect 431 -157 432 -156
rect 432 -157 433 -156
rect 433 -157 434 -156
rect 434 -157 435 -156
rect 435 -157 436 -156
rect 436 -157 437 -156
rect 437 -157 438 -156
rect 438 -157 439 -156
rect 439 -157 440 -156
rect 440 -157 441 -156
rect 441 -157 442 -156
rect 442 -157 443 -156
rect 443 -157 444 -156
rect 444 -157 445 -156
rect 445 -157 446 -156
rect 446 -157 447 -156
rect 447 -157 448 -156
rect 448 -157 449 -156
rect 449 -157 450 -156
rect 450 -157 451 -156
rect 451 -157 452 -156
rect 452 -157 453 -156
rect 453 -157 454 -156
rect 454 -157 455 -156
rect 455 -157 456 -156
rect 456 -157 457 -156
rect 457 -157 458 -156
rect 458 -157 459 -156
rect 459 -157 460 -156
rect 460 -157 461 -156
rect 461 -157 462 -156
rect 462 -157 463 -156
rect 463 -157 464 -156
rect 464 -157 465 -156
rect 465 -157 466 -156
rect 466 -157 467 -156
rect 467 -157 468 -156
rect 468 -157 469 -156
rect 469 -157 470 -156
rect 470 -157 471 -156
rect 471 -157 472 -156
rect 472 -157 473 -156
rect 473 -157 474 -156
rect 474 -157 475 -156
rect 475 -157 476 -156
rect 476 -157 477 -156
rect 477 -157 478 -156
rect 478 -157 479 -156
rect 479 -157 480 -156
rect 2 -158 3 -157
rect 3 -158 4 -157
rect 4 -158 5 -157
rect 5 -158 6 -157
rect 6 -158 7 -157
rect 7 -158 8 -157
rect 8 -158 9 -157
rect 9 -158 10 -157
rect 10 -158 11 -157
rect 11 -158 12 -157
rect 12 -158 13 -157
rect 13 -158 14 -157
rect 14 -158 15 -157
rect 15 -158 16 -157
rect 16 -158 17 -157
rect 17 -158 18 -157
rect 18 -158 19 -157
rect 19 -158 20 -157
rect 20 -158 21 -157
rect 21 -158 22 -157
rect 22 -158 23 -157
rect 23 -158 24 -157
rect 24 -158 25 -157
rect 25 -158 26 -157
rect 26 -158 27 -157
rect 27 -158 28 -157
rect 28 -158 29 -157
rect 29 -158 30 -157
rect 30 -158 31 -157
rect 31 -158 32 -157
rect 32 -158 33 -157
rect 33 -158 34 -157
rect 34 -158 35 -157
rect 35 -158 36 -157
rect 36 -158 37 -157
rect 37 -158 38 -157
rect 38 -158 39 -157
rect 39 -158 40 -157
rect 40 -158 41 -157
rect 41 -158 42 -157
rect 42 -158 43 -157
rect 43 -158 44 -157
rect 44 -158 45 -157
rect 45 -158 46 -157
rect 46 -158 47 -157
rect 47 -158 48 -157
rect 48 -158 49 -157
rect 49 -158 50 -157
rect 50 -158 51 -157
rect 51 -158 52 -157
rect 52 -158 53 -157
rect 53 -158 54 -157
rect 54 -158 55 -157
rect 55 -158 56 -157
rect 56 -158 57 -157
rect 57 -158 58 -157
rect 58 -158 59 -157
rect 59 -158 60 -157
rect 60 -158 61 -157
rect 61 -158 62 -157
rect 62 -158 63 -157
rect 63 -158 64 -157
rect 64 -158 65 -157
rect 65 -158 66 -157
rect 66 -158 67 -157
rect 67 -158 68 -157
rect 68 -158 69 -157
rect 69 -158 70 -157
rect 70 -158 71 -157
rect 71 -158 72 -157
rect 72 -158 73 -157
rect 73 -158 74 -157
rect 74 -158 75 -157
rect 75 -158 76 -157
rect 76 -158 77 -157
rect 77 -158 78 -157
rect 78 -158 79 -157
rect 79 -158 80 -157
rect 80 -158 81 -157
rect 81 -158 82 -157
rect 82 -158 83 -157
rect 83 -158 84 -157
rect 84 -158 85 -157
rect 85 -158 86 -157
rect 86 -158 87 -157
rect 87 -158 88 -157
rect 88 -158 89 -157
rect 89 -158 90 -157
rect 90 -158 91 -157
rect 91 -158 92 -157
rect 92 -158 93 -157
rect 93 -158 94 -157
rect 94 -158 95 -157
rect 95 -158 96 -157
rect 96 -158 97 -157
rect 97 -158 98 -157
rect 98 -158 99 -157
rect 99 -158 100 -157
rect 100 -158 101 -157
rect 101 -158 102 -157
rect 102 -158 103 -157
rect 103 -158 104 -157
rect 104 -158 105 -157
rect 105 -158 106 -157
rect 106 -158 107 -157
rect 107 -158 108 -157
rect 108 -158 109 -157
rect 109 -158 110 -157
rect 110 -158 111 -157
rect 111 -158 112 -157
rect 112 -158 113 -157
rect 113 -158 114 -157
rect 114 -158 115 -157
rect 115 -158 116 -157
rect 116 -158 117 -157
rect 117 -158 118 -157
rect 118 -158 119 -157
rect 119 -158 120 -157
rect 120 -158 121 -157
rect 121 -158 122 -157
rect 122 -158 123 -157
rect 123 -158 124 -157
rect 124 -158 125 -157
rect 125 -158 126 -157
rect 126 -158 127 -157
rect 127 -158 128 -157
rect 128 -158 129 -157
rect 129 -158 130 -157
rect 130 -158 131 -157
rect 131 -158 132 -157
rect 132 -158 133 -157
rect 133 -158 134 -157
rect 134 -158 135 -157
rect 135 -158 136 -157
rect 136 -158 137 -157
rect 137 -158 138 -157
rect 138 -158 139 -157
rect 139 -158 140 -157
rect 140 -158 141 -157
rect 141 -158 142 -157
rect 142 -158 143 -157
rect 143 -158 144 -157
rect 144 -158 145 -157
rect 145 -158 146 -157
rect 146 -158 147 -157
rect 147 -158 148 -157
rect 148 -158 149 -157
rect 149 -158 150 -157
rect 150 -158 151 -157
rect 151 -158 152 -157
rect 152 -158 153 -157
rect 153 -158 154 -157
rect 154 -158 155 -157
rect 155 -158 156 -157
rect 156 -158 157 -157
rect 157 -158 158 -157
rect 158 -158 159 -157
rect 159 -158 160 -157
rect 160 -158 161 -157
rect 161 -158 162 -157
rect 162 -158 163 -157
rect 163 -158 164 -157
rect 164 -158 165 -157
rect 165 -158 166 -157
rect 166 -158 167 -157
rect 167 -158 168 -157
rect 168 -158 169 -157
rect 169 -158 170 -157
rect 170 -158 171 -157
rect 171 -158 172 -157
rect 172 -158 173 -157
rect 173 -158 174 -157
rect 174 -158 175 -157
rect 175 -158 176 -157
rect 176 -158 177 -157
rect 177 -158 178 -157
rect 178 -158 179 -157
rect 179 -158 180 -157
rect 180 -158 181 -157
rect 181 -158 182 -157
rect 182 -158 183 -157
rect 183 -158 184 -157
rect 184 -158 185 -157
rect 185 -158 186 -157
rect 186 -158 187 -157
rect 187 -158 188 -157
rect 188 -158 189 -157
rect 189 -158 190 -157
rect 190 -158 191 -157
rect 191 -158 192 -157
rect 192 -158 193 -157
rect 193 -158 194 -157
rect 194 -158 195 -157
rect 195 -158 196 -157
rect 196 -158 197 -157
rect 197 -158 198 -157
rect 198 -158 199 -157
rect 199 -158 200 -157
rect 200 -158 201 -157
rect 201 -158 202 -157
rect 202 -158 203 -157
rect 203 -158 204 -157
rect 204 -158 205 -157
rect 205 -158 206 -157
rect 206 -158 207 -157
rect 207 -158 208 -157
rect 208 -158 209 -157
rect 209 -158 210 -157
rect 210 -158 211 -157
rect 211 -158 212 -157
rect 212 -158 213 -157
rect 213 -158 214 -157
rect 214 -158 215 -157
rect 215 -158 216 -157
rect 216 -158 217 -157
rect 217 -158 218 -157
rect 218 -158 219 -157
rect 219 -158 220 -157
rect 220 -158 221 -157
rect 221 -158 222 -157
rect 222 -158 223 -157
rect 223 -158 224 -157
rect 224 -158 225 -157
rect 225 -158 226 -157
rect 226 -158 227 -157
rect 227 -158 228 -157
rect 228 -158 229 -157
rect 229 -158 230 -157
rect 230 -158 231 -157
rect 231 -158 232 -157
rect 232 -158 233 -157
rect 233 -158 234 -157
rect 234 -158 235 -157
rect 235 -158 236 -157
rect 236 -158 237 -157
rect 237 -158 238 -157
rect 238 -158 239 -157
rect 239 -158 240 -157
rect 240 -158 241 -157
rect 241 -158 242 -157
rect 242 -158 243 -157
rect 243 -158 244 -157
rect 244 -158 245 -157
rect 245 -158 246 -157
rect 246 -158 247 -157
rect 247 -158 248 -157
rect 248 -158 249 -157
rect 249 -158 250 -157
rect 250 -158 251 -157
rect 251 -158 252 -157
rect 252 -158 253 -157
rect 253 -158 254 -157
rect 254 -158 255 -157
rect 255 -158 256 -157
rect 256 -158 257 -157
rect 257 -158 258 -157
rect 258 -158 259 -157
rect 259 -158 260 -157
rect 260 -158 261 -157
rect 261 -158 262 -157
rect 262 -158 263 -157
rect 263 -158 264 -157
rect 264 -158 265 -157
rect 265 -158 266 -157
rect 266 -158 267 -157
rect 267 -158 268 -157
rect 268 -158 269 -157
rect 269 -158 270 -157
rect 270 -158 271 -157
rect 271 -158 272 -157
rect 272 -158 273 -157
rect 273 -158 274 -157
rect 274 -158 275 -157
rect 275 -158 276 -157
rect 276 -158 277 -157
rect 277 -158 278 -157
rect 278 -158 279 -157
rect 279 -158 280 -157
rect 280 -158 281 -157
rect 281 -158 282 -157
rect 282 -158 283 -157
rect 283 -158 284 -157
rect 284 -158 285 -157
rect 285 -158 286 -157
rect 286 -158 287 -157
rect 287 -158 288 -157
rect 288 -158 289 -157
rect 289 -158 290 -157
rect 290 -158 291 -157
rect 291 -158 292 -157
rect 292 -158 293 -157
rect 293 -158 294 -157
rect 294 -158 295 -157
rect 295 -158 296 -157
rect 296 -158 297 -157
rect 297 -158 298 -157
rect 298 -158 299 -157
rect 299 -158 300 -157
rect 300 -158 301 -157
rect 301 -158 302 -157
rect 302 -158 303 -157
rect 303 -158 304 -157
rect 304 -158 305 -157
rect 305 -158 306 -157
rect 306 -158 307 -157
rect 307 -158 308 -157
rect 308 -158 309 -157
rect 309 -158 310 -157
rect 310 -158 311 -157
rect 311 -158 312 -157
rect 312 -158 313 -157
rect 313 -158 314 -157
rect 314 -158 315 -157
rect 315 -158 316 -157
rect 316 -158 317 -157
rect 317 -158 318 -157
rect 318 -158 319 -157
rect 319 -158 320 -157
rect 320 -158 321 -157
rect 321 -158 322 -157
rect 322 -158 323 -157
rect 323 -158 324 -157
rect 324 -158 325 -157
rect 325 -158 326 -157
rect 326 -158 327 -157
rect 327 -158 328 -157
rect 328 -158 329 -157
rect 329 -158 330 -157
rect 330 -158 331 -157
rect 331 -158 332 -157
rect 332 -158 333 -157
rect 333 -158 334 -157
rect 334 -158 335 -157
rect 335 -158 336 -157
rect 336 -158 337 -157
rect 337 -158 338 -157
rect 338 -158 339 -157
rect 339 -158 340 -157
rect 340 -158 341 -157
rect 341 -158 342 -157
rect 342 -158 343 -157
rect 343 -158 344 -157
rect 344 -158 345 -157
rect 345 -158 346 -157
rect 346 -158 347 -157
rect 347 -158 348 -157
rect 348 -158 349 -157
rect 349 -158 350 -157
rect 350 -158 351 -157
rect 351 -158 352 -157
rect 352 -158 353 -157
rect 353 -158 354 -157
rect 354 -158 355 -157
rect 355 -158 356 -157
rect 356 -158 357 -157
rect 357 -158 358 -157
rect 358 -158 359 -157
rect 359 -158 360 -157
rect 360 -158 361 -157
rect 361 -158 362 -157
rect 362 -158 363 -157
rect 363 -158 364 -157
rect 364 -158 365 -157
rect 365 -158 366 -157
rect 366 -158 367 -157
rect 367 -158 368 -157
rect 368 -158 369 -157
rect 369 -158 370 -157
rect 370 -158 371 -157
rect 371 -158 372 -157
rect 372 -158 373 -157
rect 373 -158 374 -157
rect 374 -158 375 -157
rect 375 -158 376 -157
rect 376 -158 377 -157
rect 377 -158 378 -157
rect 378 -158 379 -157
rect 379 -158 380 -157
rect 380 -158 381 -157
rect 381 -158 382 -157
rect 382 -158 383 -157
rect 383 -158 384 -157
rect 384 -158 385 -157
rect 385 -158 386 -157
rect 386 -158 387 -157
rect 387 -158 388 -157
rect 388 -158 389 -157
rect 389 -158 390 -157
rect 390 -158 391 -157
rect 391 -158 392 -157
rect 392 -158 393 -157
rect 393 -158 394 -157
rect 394 -158 395 -157
rect 395 -158 396 -157
rect 396 -158 397 -157
rect 397 -158 398 -157
rect 398 -158 399 -157
rect 399 -158 400 -157
rect 400 -158 401 -157
rect 401 -158 402 -157
rect 402 -158 403 -157
rect 403 -158 404 -157
rect 404 -158 405 -157
rect 405 -158 406 -157
rect 406 -158 407 -157
rect 407 -158 408 -157
rect 408 -158 409 -157
rect 409 -158 410 -157
rect 410 -158 411 -157
rect 411 -158 412 -157
rect 412 -158 413 -157
rect 413 -158 414 -157
rect 414 -158 415 -157
rect 415 -158 416 -157
rect 416 -158 417 -157
rect 417 -158 418 -157
rect 418 -158 419 -157
rect 419 -158 420 -157
rect 420 -158 421 -157
rect 421 -158 422 -157
rect 422 -158 423 -157
rect 423 -158 424 -157
rect 424 -158 425 -157
rect 425 -158 426 -157
rect 426 -158 427 -157
rect 427 -158 428 -157
rect 428 -158 429 -157
rect 429 -158 430 -157
rect 430 -158 431 -157
rect 431 -158 432 -157
rect 432 -158 433 -157
rect 433 -158 434 -157
rect 434 -158 435 -157
rect 435 -158 436 -157
rect 436 -158 437 -157
rect 437 -158 438 -157
rect 438 -158 439 -157
rect 439 -158 440 -157
rect 440 -158 441 -157
rect 441 -158 442 -157
rect 442 -158 443 -157
rect 443 -158 444 -157
rect 444 -158 445 -157
rect 445 -158 446 -157
rect 446 -158 447 -157
rect 447 -158 448 -157
rect 448 -158 449 -157
rect 449 -158 450 -157
rect 450 -158 451 -157
rect 451 -158 452 -157
rect 452 -158 453 -157
rect 453 -158 454 -157
rect 454 -158 455 -157
rect 455 -158 456 -157
rect 456 -158 457 -157
rect 457 -158 458 -157
rect 458 -158 459 -157
rect 459 -158 460 -157
rect 460 -158 461 -157
rect 461 -158 462 -157
rect 462 -158 463 -157
rect 463 -158 464 -157
rect 464 -158 465 -157
rect 465 -158 466 -157
rect 466 -158 467 -157
rect 467 -158 468 -157
rect 468 -158 469 -157
rect 469 -158 470 -157
rect 470 -158 471 -157
rect 471 -158 472 -157
rect 472 -158 473 -157
rect 473 -158 474 -157
rect 474 -158 475 -157
rect 475 -158 476 -157
rect 476 -158 477 -157
rect 477 -158 478 -157
rect 478 -158 479 -157
rect 479 -158 480 -157
rect 2 -159 3 -158
rect 3 -159 4 -158
rect 4 -159 5 -158
rect 5 -159 6 -158
rect 6 -159 7 -158
rect 7 -159 8 -158
rect 8 -159 9 -158
rect 9 -159 10 -158
rect 10 -159 11 -158
rect 11 -159 12 -158
rect 12 -159 13 -158
rect 13 -159 14 -158
rect 14 -159 15 -158
rect 15 -159 16 -158
rect 16 -159 17 -158
rect 17 -159 18 -158
rect 18 -159 19 -158
rect 19 -159 20 -158
rect 20 -159 21 -158
rect 21 -159 22 -158
rect 22 -159 23 -158
rect 23 -159 24 -158
rect 24 -159 25 -158
rect 25 -159 26 -158
rect 26 -159 27 -158
rect 27 -159 28 -158
rect 28 -159 29 -158
rect 29 -159 30 -158
rect 30 -159 31 -158
rect 31 -159 32 -158
rect 32 -159 33 -158
rect 33 -159 34 -158
rect 34 -159 35 -158
rect 35 -159 36 -158
rect 36 -159 37 -158
rect 37 -159 38 -158
rect 38 -159 39 -158
rect 39 -159 40 -158
rect 40 -159 41 -158
rect 41 -159 42 -158
rect 42 -159 43 -158
rect 43 -159 44 -158
rect 44 -159 45 -158
rect 45 -159 46 -158
rect 46 -159 47 -158
rect 47 -159 48 -158
rect 48 -159 49 -158
rect 49 -159 50 -158
rect 50 -159 51 -158
rect 51 -159 52 -158
rect 52 -159 53 -158
rect 53 -159 54 -158
rect 54 -159 55 -158
rect 55 -159 56 -158
rect 56 -159 57 -158
rect 57 -159 58 -158
rect 58 -159 59 -158
rect 59 -159 60 -158
rect 60 -159 61 -158
rect 61 -159 62 -158
rect 62 -159 63 -158
rect 63 -159 64 -158
rect 64 -159 65 -158
rect 65 -159 66 -158
rect 66 -159 67 -158
rect 67 -159 68 -158
rect 68 -159 69 -158
rect 69 -159 70 -158
rect 70 -159 71 -158
rect 71 -159 72 -158
rect 72 -159 73 -158
rect 73 -159 74 -158
rect 74 -159 75 -158
rect 75 -159 76 -158
rect 76 -159 77 -158
rect 77 -159 78 -158
rect 78 -159 79 -158
rect 79 -159 80 -158
rect 80 -159 81 -158
rect 81 -159 82 -158
rect 82 -159 83 -158
rect 83 -159 84 -158
rect 84 -159 85 -158
rect 85 -159 86 -158
rect 86 -159 87 -158
rect 87 -159 88 -158
rect 88 -159 89 -158
rect 89 -159 90 -158
rect 90 -159 91 -158
rect 91 -159 92 -158
rect 92 -159 93 -158
rect 93 -159 94 -158
rect 94 -159 95 -158
rect 95 -159 96 -158
rect 96 -159 97 -158
rect 97 -159 98 -158
rect 98 -159 99 -158
rect 99 -159 100 -158
rect 100 -159 101 -158
rect 101 -159 102 -158
rect 102 -159 103 -158
rect 103 -159 104 -158
rect 104 -159 105 -158
rect 105 -159 106 -158
rect 106 -159 107 -158
rect 107 -159 108 -158
rect 108 -159 109 -158
rect 109 -159 110 -158
rect 110 -159 111 -158
rect 111 -159 112 -158
rect 112 -159 113 -158
rect 113 -159 114 -158
rect 114 -159 115 -158
rect 115 -159 116 -158
rect 116 -159 117 -158
rect 117 -159 118 -158
rect 118 -159 119 -158
rect 119 -159 120 -158
rect 120 -159 121 -158
rect 121 -159 122 -158
rect 122 -159 123 -158
rect 123 -159 124 -158
rect 124 -159 125 -158
rect 125 -159 126 -158
rect 126 -159 127 -158
rect 127 -159 128 -158
rect 128 -159 129 -158
rect 129 -159 130 -158
rect 130 -159 131 -158
rect 131 -159 132 -158
rect 132 -159 133 -158
rect 133 -159 134 -158
rect 134 -159 135 -158
rect 135 -159 136 -158
rect 136 -159 137 -158
rect 137 -159 138 -158
rect 138 -159 139 -158
rect 139 -159 140 -158
rect 140 -159 141 -158
rect 141 -159 142 -158
rect 142 -159 143 -158
rect 143 -159 144 -158
rect 144 -159 145 -158
rect 145 -159 146 -158
rect 146 -159 147 -158
rect 147 -159 148 -158
rect 148 -159 149 -158
rect 149 -159 150 -158
rect 150 -159 151 -158
rect 151 -159 152 -158
rect 152 -159 153 -158
rect 153 -159 154 -158
rect 154 -159 155 -158
rect 155 -159 156 -158
rect 156 -159 157 -158
rect 157 -159 158 -158
rect 158 -159 159 -158
rect 159 -159 160 -158
rect 160 -159 161 -158
rect 161 -159 162 -158
rect 162 -159 163 -158
rect 163 -159 164 -158
rect 164 -159 165 -158
rect 165 -159 166 -158
rect 166 -159 167 -158
rect 167 -159 168 -158
rect 168 -159 169 -158
rect 169 -159 170 -158
rect 170 -159 171 -158
rect 171 -159 172 -158
rect 172 -159 173 -158
rect 173 -159 174 -158
rect 174 -159 175 -158
rect 175 -159 176 -158
rect 176 -159 177 -158
rect 177 -159 178 -158
rect 178 -159 179 -158
rect 179 -159 180 -158
rect 180 -159 181 -158
rect 181 -159 182 -158
rect 182 -159 183 -158
rect 183 -159 184 -158
rect 184 -159 185 -158
rect 185 -159 186 -158
rect 186 -159 187 -158
rect 187 -159 188 -158
rect 188 -159 189 -158
rect 189 -159 190 -158
rect 190 -159 191 -158
rect 191 -159 192 -158
rect 192 -159 193 -158
rect 193 -159 194 -158
rect 194 -159 195 -158
rect 195 -159 196 -158
rect 196 -159 197 -158
rect 197 -159 198 -158
rect 198 -159 199 -158
rect 199 -159 200 -158
rect 200 -159 201 -158
rect 201 -159 202 -158
rect 202 -159 203 -158
rect 203 -159 204 -158
rect 204 -159 205 -158
rect 205 -159 206 -158
rect 206 -159 207 -158
rect 207 -159 208 -158
rect 208 -159 209 -158
rect 209 -159 210 -158
rect 210 -159 211 -158
rect 211 -159 212 -158
rect 212 -159 213 -158
rect 213 -159 214 -158
rect 214 -159 215 -158
rect 215 -159 216 -158
rect 216 -159 217 -158
rect 217 -159 218 -158
rect 218 -159 219 -158
rect 219 -159 220 -158
rect 220 -159 221 -158
rect 221 -159 222 -158
rect 222 -159 223 -158
rect 223 -159 224 -158
rect 224 -159 225 -158
rect 225 -159 226 -158
rect 226 -159 227 -158
rect 227 -159 228 -158
rect 228 -159 229 -158
rect 229 -159 230 -158
rect 230 -159 231 -158
rect 231 -159 232 -158
rect 232 -159 233 -158
rect 233 -159 234 -158
rect 234 -159 235 -158
rect 235 -159 236 -158
rect 236 -159 237 -158
rect 237 -159 238 -158
rect 238 -159 239 -158
rect 239 -159 240 -158
rect 240 -159 241 -158
rect 241 -159 242 -158
rect 242 -159 243 -158
rect 243 -159 244 -158
rect 244 -159 245 -158
rect 245 -159 246 -158
rect 246 -159 247 -158
rect 247 -159 248 -158
rect 248 -159 249 -158
rect 249 -159 250 -158
rect 250 -159 251 -158
rect 251 -159 252 -158
rect 252 -159 253 -158
rect 253 -159 254 -158
rect 254 -159 255 -158
rect 255 -159 256 -158
rect 256 -159 257 -158
rect 257 -159 258 -158
rect 258 -159 259 -158
rect 259 -159 260 -158
rect 260 -159 261 -158
rect 261 -159 262 -158
rect 262 -159 263 -158
rect 263 -159 264 -158
rect 264 -159 265 -158
rect 265 -159 266 -158
rect 266 -159 267 -158
rect 267 -159 268 -158
rect 268 -159 269 -158
rect 269 -159 270 -158
rect 270 -159 271 -158
rect 271 -159 272 -158
rect 272 -159 273 -158
rect 273 -159 274 -158
rect 274 -159 275 -158
rect 275 -159 276 -158
rect 276 -159 277 -158
rect 277 -159 278 -158
rect 278 -159 279 -158
rect 279 -159 280 -158
rect 280 -159 281 -158
rect 281 -159 282 -158
rect 282 -159 283 -158
rect 283 -159 284 -158
rect 284 -159 285 -158
rect 285 -159 286 -158
rect 286 -159 287 -158
rect 287 -159 288 -158
rect 288 -159 289 -158
rect 289 -159 290 -158
rect 290 -159 291 -158
rect 291 -159 292 -158
rect 292 -159 293 -158
rect 293 -159 294 -158
rect 294 -159 295 -158
rect 295 -159 296 -158
rect 296 -159 297 -158
rect 297 -159 298 -158
rect 298 -159 299 -158
rect 299 -159 300 -158
rect 300 -159 301 -158
rect 301 -159 302 -158
rect 302 -159 303 -158
rect 303 -159 304 -158
rect 304 -159 305 -158
rect 305 -159 306 -158
rect 306 -159 307 -158
rect 307 -159 308 -158
rect 308 -159 309 -158
rect 309 -159 310 -158
rect 310 -159 311 -158
rect 311 -159 312 -158
rect 312 -159 313 -158
rect 313 -159 314 -158
rect 314 -159 315 -158
rect 315 -159 316 -158
rect 316 -159 317 -158
rect 317 -159 318 -158
rect 318 -159 319 -158
rect 319 -159 320 -158
rect 320 -159 321 -158
rect 321 -159 322 -158
rect 322 -159 323 -158
rect 323 -159 324 -158
rect 324 -159 325 -158
rect 325 -159 326 -158
rect 326 -159 327 -158
rect 327 -159 328 -158
rect 328 -159 329 -158
rect 329 -159 330 -158
rect 330 -159 331 -158
rect 331 -159 332 -158
rect 332 -159 333 -158
rect 333 -159 334 -158
rect 334 -159 335 -158
rect 335 -159 336 -158
rect 336 -159 337 -158
rect 337 -159 338 -158
rect 338 -159 339 -158
rect 339 -159 340 -158
rect 340 -159 341 -158
rect 341 -159 342 -158
rect 342 -159 343 -158
rect 343 -159 344 -158
rect 344 -159 345 -158
rect 345 -159 346 -158
rect 346 -159 347 -158
rect 347 -159 348 -158
rect 348 -159 349 -158
rect 349 -159 350 -158
rect 350 -159 351 -158
rect 351 -159 352 -158
rect 352 -159 353 -158
rect 353 -159 354 -158
rect 354 -159 355 -158
rect 355 -159 356 -158
rect 356 -159 357 -158
rect 357 -159 358 -158
rect 358 -159 359 -158
rect 359 -159 360 -158
rect 360 -159 361 -158
rect 361 -159 362 -158
rect 362 -159 363 -158
rect 363 -159 364 -158
rect 364 -159 365 -158
rect 365 -159 366 -158
rect 366 -159 367 -158
rect 367 -159 368 -158
rect 368 -159 369 -158
rect 369 -159 370 -158
rect 370 -159 371 -158
rect 371 -159 372 -158
rect 372 -159 373 -158
rect 373 -159 374 -158
rect 374 -159 375 -158
rect 375 -159 376 -158
rect 376 -159 377 -158
rect 377 -159 378 -158
rect 378 -159 379 -158
rect 379 -159 380 -158
rect 380 -159 381 -158
rect 381 -159 382 -158
rect 382 -159 383 -158
rect 383 -159 384 -158
rect 384 -159 385 -158
rect 385 -159 386 -158
rect 386 -159 387 -158
rect 387 -159 388 -158
rect 388 -159 389 -158
rect 389 -159 390 -158
rect 390 -159 391 -158
rect 391 -159 392 -158
rect 392 -159 393 -158
rect 393 -159 394 -158
rect 394 -159 395 -158
rect 395 -159 396 -158
rect 396 -159 397 -158
rect 397 -159 398 -158
rect 398 -159 399 -158
rect 399 -159 400 -158
rect 400 -159 401 -158
rect 401 -159 402 -158
rect 402 -159 403 -158
rect 403 -159 404 -158
rect 404 -159 405 -158
rect 405 -159 406 -158
rect 406 -159 407 -158
rect 407 -159 408 -158
rect 408 -159 409 -158
rect 409 -159 410 -158
rect 410 -159 411 -158
rect 411 -159 412 -158
rect 412 -159 413 -158
rect 413 -159 414 -158
rect 414 -159 415 -158
rect 415 -159 416 -158
rect 416 -159 417 -158
rect 417 -159 418 -158
rect 418 -159 419 -158
rect 419 -159 420 -158
rect 420 -159 421 -158
rect 421 -159 422 -158
rect 422 -159 423 -158
rect 423 -159 424 -158
rect 424 -159 425 -158
rect 425 -159 426 -158
rect 426 -159 427 -158
rect 427 -159 428 -158
rect 428 -159 429 -158
rect 429 -159 430 -158
rect 430 -159 431 -158
rect 431 -159 432 -158
rect 432 -159 433 -158
rect 433 -159 434 -158
rect 434 -159 435 -158
rect 435 -159 436 -158
rect 436 -159 437 -158
rect 437 -159 438 -158
rect 438 -159 439 -158
rect 439 -159 440 -158
rect 440 -159 441 -158
rect 441 -159 442 -158
rect 442 -159 443 -158
rect 443 -159 444 -158
rect 444 -159 445 -158
rect 445 -159 446 -158
rect 446 -159 447 -158
rect 447 -159 448 -158
rect 448 -159 449 -158
rect 449 -159 450 -158
rect 450 -159 451 -158
rect 451 -159 452 -158
rect 452 -159 453 -158
rect 453 -159 454 -158
rect 454 -159 455 -158
rect 455 -159 456 -158
rect 456 -159 457 -158
rect 457 -159 458 -158
rect 458 -159 459 -158
rect 459 -159 460 -158
rect 460 -159 461 -158
rect 461 -159 462 -158
rect 462 -159 463 -158
rect 463 -159 464 -158
rect 464 -159 465 -158
rect 465 -159 466 -158
rect 466 -159 467 -158
rect 467 -159 468 -158
rect 468 -159 469 -158
rect 469 -159 470 -158
rect 470 -159 471 -158
rect 471 -159 472 -158
rect 472 -159 473 -158
rect 473 -159 474 -158
rect 474 -159 475 -158
rect 475 -159 476 -158
rect 476 -159 477 -158
rect 477 -159 478 -158
rect 478 -159 479 -158
rect 479 -159 480 -158
rect 2 -160 3 -159
rect 3 -160 4 -159
rect 4 -160 5 -159
rect 5 -160 6 -159
rect 6 -160 7 -159
rect 7 -160 8 -159
rect 8 -160 9 -159
rect 9 -160 10 -159
rect 10 -160 11 -159
rect 11 -160 12 -159
rect 12 -160 13 -159
rect 13 -160 14 -159
rect 14 -160 15 -159
rect 15 -160 16 -159
rect 16 -160 17 -159
rect 17 -160 18 -159
rect 18 -160 19 -159
rect 19 -160 20 -159
rect 20 -160 21 -159
rect 21 -160 22 -159
rect 22 -160 23 -159
rect 23 -160 24 -159
rect 24 -160 25 -159
rect 25 -160 26 -159
rect 26 -160 27 -159
rect 27 -160 28 -159
rect 28 -160 29 -159
rect 29 -160 30 -159
rect 30 -160 31 -159
rect 31 -160 32 -159
rect 32 -160 33 -159
rect 33 -160 34 -159
rect 34 -160 35 -159
rect 35 -160 36 -159
rect 36 -160 37 -159
rect 37 -160 38 -159
rect 38 -160 39 -159
rect 39 -160 40 -159
rect 40 -160 41 -159
rect 41 -160 42 -159
rect 42 -160 43 -159
rect 43 -160 44 -159
rect 44 -160 45 -159
rect 45 -160 46 -159
rect 46 -160 47 -159
rect 47 -160 48 -159
rect 48 -160 49 -159
rect 49 -160 50 -159
rect 50 -160 51 -159
rect 51 -160 52 -159
rect 52 -160 53 -159
rect 53 -160 54 -159
rect 54 -160 55 -159
rect 55 -160 56 -159
rect 56 -160 57 -159
rect 57 -160 58 -159
rect 58 -160 59 -159
rect 59 -160 60 -159
rect 60 -160 61 -159
rect 61 -160 62 -159
rect 62 -160 63 -159
rect 63 -160 64 -159
rect 64 -160 65 -159
rect 65 -160 66 -159
rect 66 -160 67 -159
rect 67 -160 68 -159
rect 68 -160 69 -159
rect 69 -160 70 -159
rect 70 -160 71 -159
rect 71 -160 72 -159
rect 72 -160 73 -159
rect 73 -160 74 -159
rect 74 -160 75 -159
rect 75 -160 76 -159
rect 76 -160 77 -159
rect 77 -160 78 -159
rect 78 -160 79 -159
rect 79 -160 80 -159
rect 80 -160 81 -159
rect 81 -160 82 -159
rect 82 -160 83 -159
rect 83 -160 84 -159
rect 84 -160 85 -159
rect 85 -160 86 -159
rect 86 -160 87 -159
rect 87 -160 88 -159
rect 88 -160 89 -159
rect 89 -160 90 -159
rect 90 -160 91 -159
rect 91 -160 92 -159
rect 92 -160 93 -159
rect 93 -160 94 -159
rect 94 -160 95 -159
rect 95 -160 96 -159
rect 96 -160 97 -159
rect 97 -160 98 -159
rect 98 -160 99 -159
rect 99 -160 100 -159
rect 100 -160 101 -159
rect 101 -160 102 -159
rect 102 -160 103 -159
rect 103 -160 104 -159
rect 104 -160 105 -159
rect 105 -160 106 -159
rect 106 -160 107 -159
rect 107 -160 108 -159
rect 108 -160 109 -159
rect 109 -160 110 -159
rect 110 -160 111 -159
rect 111 -160 112 -159
rect 112 -160 113 -159
rect 113 -160 114 -159
rect 114 -160 115 -159
rect 115 -160 116 -159
rect 116 -160 117 -159
rect 117 -160 118 -159
rect 118 -160 119 -159
rect 119 -160 120 -159
rect 120 -160 121 -159
rect 121 -160 122 -159
rect 122 -160 123 -159
rect 123 -160 124 -159
rect 124 -160 125 -159
rect 125 -160 126 -159
rect 126 -160 127 -159
rect 127 -160 128 -159
rect 128 -160 129 -159
rect 129 -160 130 -159
rect 130 -160 131 -159
rect 131 -160 132 -159
rect 132 -160 133 -159
rect 133 -160 134 -159
rect 134 -160 135 -159
rect 135 -160 136 -159
rect 136 -160 137 -159
rect 137 -160 138 -159
rect 138 -160 139 -159
rect 139 -160 140 -159
rect 140 -160 141 -159
rect 141 -160 142 -159
rect 142 -160 143 -159
rect 143 -160 144 -159
rect 144 -160 145 -159
rect 145 -160 146 -159
rect 146 -160 147 -159
rect 147 -160 148 -159
rect 148 -160 149 -159
rect 149 -160 150 -159
rect 150 -160 151 -159
rect 151 -160 152 -159
rect 152 -160 153 -159
rect 153 -160 154 -159
rect 154 -160 155 -159
rect 155 -160 156 -159
rect 156 -160 157 -159
rect 157 -160 158 -159
rect 158 -160 159 -159
rect 159 -160 160 -159
rect 160 -160 161 -159
rect 161 -160 162 -159
rect 162 -160 163 -159
rect 163 -160 164 -159
rect 164 -160 165 -159
rect 165 -160 166 -159
rect 166 -160 167 -159
rect 167 -160 168 -159
rect 168 -160 169 -159
rect 169 -160 170 -159
rect 170 -160 171 -159
rect 171 -160 172 -159
rect 172 -160 173 -159
rect 173 -160 174 -159
rect 174 -160 175 -159
rect 175 -160 176 -159
rect 176 -160 177 -159
rect 177 -160 178 -159
rect 178 -160 179 -159
rect 179 -160 180 -159
rect 180 -160 181 -159
rect 181 -160 182 -159
rect 182 -160 183 -159
rect 183 -160 184 -159
rect 184 -160 185 -159
rect 185 -160 186 -159
rect 186 -160 187 -159
rect 187 -160 188 -159
rect 188 -160 189 -159
rect 189 -160 190 -159
rect 190 -160 191 -159
rect 191 -160 192 -159
rect 192 -160 193 -159
rect 193 -160 194 -159
rect 194 -160 195 -159
rect 195 -160 196 -159
rect 196 -160 197 -159
rect 197 -160 198 -159
rect 198 -160 199 -159
rect 199 -160 200 -159
rect 200 -160 201 -159
rect 201 -160 202 -159
rect 202 -160 203 -159
rect 203 -160 204 -159
rect 204 -160 205 -159
rect 205 -160 206 -159
rect 206 -160 207 -159
rect 207 -160 208 -159
rect 208 -160 209 -159
rect 209 -160 210 -159
rect 210 -160 211 -159
rect 211 -160 212 -159
rect 212 -160 213 -159
rect 213 -160 214 -159
rect 214 -160 215 -159
rect 215 -160 216 -159
rect 216 -160 217 -159
rect 217 -160 218 -159
rect 218 -160 219 -159
rect 219 -160 220 -159
rect 220 -160 221 -159
rect 221 -160 222 -159
rect 222 -160 223 -159
rect 223 -160 224 -159
rect 224 -160 225 -159
rect 225 -160 226 -159
rect 226 -160 227 -159
rect 227 -160 228 -159
rect 228 -160 229 -159
rect 229 -160 230 -159
rect 230 -160 231 -159
rect 231 -160 232 -159
rect 232 -160 233 -159
rect 233 -160 234 -159
rect 234 -160 235 -159
rect 235 -160 236 -159
rect 236 -160 237 -159
rect 237 -160 238 -159
rect 238 -160 239 -159
rect 239 -160 240 -159
rect 240 -160 241 -159
rect 241 -160 242 -159
rect 242 -160 243 -159
rect 243 -160 244 -159
rect 244 -160 245 -159
rect 245 -160 246 -159
rect 246 -160 247 -159
rect 247 -160 248 -159
rect 248 -160 249 -159
rect 249 -160 250 -159
rect 250 -160 251 -159
rect 251 -160 252 -159
rect 252 -160 253 -159
rect 253 -160 254 -159
rect 254 -160 255 -159
rect 255 -160 256 -159
rect 256 -160 257 -159
rect 257 -160 258 -159
rect 258 -160 259 -159
rect 259 -160 260 -159
rect 260 -160 261 -159
rect 261 -160 262 -159
rect 262 -160 263 -159
rect 263 -160 264 -159
rect 264 -160 265 -159
rect 265 -160 266 -159
rect 266 -160 267 -159
rect 267 -160 268 -159
rect 268 -160 269 -159
rect 269 -160 270 -159
rect 270 -160 271 -159
rect 271 -160 272 -159
rect 272 -160 273 -159
rect 273 -160 274 -159
rect 274 -160 275 -159
rect 275 -160 276 -159
rect 276 -160 277 -159
rect 277 -160 278 -159
rect 278 -160 279 -159
rect 279 -160 280 -159
rect 280 -160 281 -159
rect 281 -160 282 -159
rect 282 -160 283 -159
rect 283 -160 284 -159
rect 284 -160 285 -159
rect 285 -160 286 -159
rect 286 -160 287 -159
rect 287 -160 288 -159
rect 288 -160 289 -159
rect 289 -160 290 -159
rect 290 -160 291 -159
rect 291 -160 292 -159
rect 292 -160 293 -159
rect 293 -160 294 -159
rect 294 -160 295 -159
rect 295 -160 296 -159
rect 296 -160 297 -159
rect 297 -160 298 -159
rect 298 -160 299 -159
rect 299 -160 300 -159
rect 300 -160 301 -159
rect 301 -160 302 -159
rect 302 -160 303 -159
rect 303 -160 304 -159
rect 304 -160 305 -159
rect 305 -160 306 -159
rect 306 -160 307 -159
rect 307 -160 308 -159
rect 308 -160 309 -159
rect 309 -160 310 -159
rect 310 -160 311 -159
rect 311 -160 312 -159
rect 312 -160 313 -159
rect 313 -160 314 -159
rect 314 -160 315 -159
rect 315 -160 316 -159
rect 316 -160 317 -159
rect 317 -160 318 -159
rect 318 -160 319 -159
rect 319 -160 320 -159
rect 320 -160 321 -159
rect 321 -160 322 -159
rect 322 -160 323 -159
rect 323 -160 324 -159
rect 324 -160 325 -159
rect 325 -160 326 -159
rect 326 -160 327 -159
rect 327 -160 328 -159
rect 328 -160 329 -159
rect 329 -160 330 -159
rect 330 -160 331 -159
rect 331 -160 332 -159
rect 332 -160 333 -159
rect 333 -160 334 -159
rect 334 -160 335 -159
rect 335 -160 336 -159
rect 336 -160 337 -159
rect 337 -160 338 -159
rect 338 -160 339 -159
rect 339 -160 340 -159
rect 340 -160 341 -159
rect 341 -160 342 -159
rect 342 -160 343 -159
rect 343 -160 344 -159
rect 344 -160 345 -159
rect 345 -160 346 -159
rect 346 -160 347 -159
rect 347 -160 348 -159
rect 348 -160 349 -159
rect 349 -160 350 -159
rect 350 -160 351 -159
rect 351 -160 352 -159
rect 352 -160 353 -159
rect 353 -160 354 -159
rect 354 -160 355 -159
rect 355 -160 356 -159
rect 356 -160 357 -159
rect 357 -160 358 -159
rect 358 -160 359 -159
rect 359 -160 360 -159
rect 360 -160 361 -159
rect 361 -160 362 -159
rect 362 -160 363 -159
rect 363 -160 364 -159
rect 364 -160 365 -159
rect 365 -160 366 -159
rect 366 -160 367 -159
rect 367 -160 368 -159
rect 368 -160 369 -159
rect 369 -160 370 -159
rect 370 -160 371 -159
rect 371 -160 372 -159
rect 372 -160 373 -159
rect 373 -160 374 -159
rect 374 -160 375 -159
rect 375 -160 376 -159
rect 376 -160 377 -159
rect 377 -160 378 -159
rect 378 -160 379 -159
rect 379 -160 380 -159
rect 380 -160 381 -159
rect 381 -160 382 -159
rect 382 -160 383 -159
rect 383 -160 384 -159
rect 384 -160 385 -159
rect 385 -160 386 -159
rect 386 -160 387 -159
rect 387 -160 388 -159
rect 388 -160 389 -159
rect 389 -160 390 -159
rect 390 -160 391 -159
rect 391 -160 392 -159
rect 392 -160 393 -159
rect 393 -160 394 -159
rect 394 -160 395 -159
rect 395 -160 396 -159
rect 396 -160 397 -159
rect 397 -160 398 -159
rect 398 -160 399 -159
rect 399 -160 400 -159
rect 400 -160 401 -159
rect 401 -160 402 -159
rect 402 -160 403 -159
rect 403 -160 404 -159
rect 404 -160 405 -159
rect 405 -160 406 -159
rect 406 -160 407 -159
rect 407 -160 408 -159
rect 408 -160 409 -159
rect 409 -160 410 -159
rect 410 -160 411 -159
rect 411 -160 412 -159
rect 412 -160 413 -159
rect 413 -160 414 -159
rect 414 -160 415 -159
rect 415 -160 416 -159
rect 416 -160 417 -159
rect 417 -160 418 -159
rect 418 -160 419 -159
rect 419 -160 420 -159
rect 420 -160 421 -159
rect 421 -160 422 -159
rect 422 -160 423 -159
rect 423 -160 424 -159
rect 424 -160 425 -159
rect 425 -160 426 -159
rect 426 -160 427 -159
rect 427 -160 428 -159
rect 428 -160 429 -159
rect 429 -160 430 -159
rect 430 -160 431 -159
rect 431 -160 432 -159
rect 432 -160 433 -159
rect 433 -160 434 -159
rect 434 -160 435 -159
rect 435 -160 436 -159
rect 436 -160 437 -159
rect 437 -160 438 -159
rect 438 -160 439 -159
rect 439 -160 440 -159
rect 440 -160 441 -159
rect 441 -160 442 -159
rect 442 -160 443 -159
rect 443 -160 444 -159
rect 444 -160 445 -159
rect 445 -160 446 -159
rect 446 -160 447 -159
rect 447 -160 448 -159
rect 448 -160 449 -159
rect 449 -160 450 -159
rect 450 -160 451 -159
rect 451 -160 452 -159
rect 452 -160 453 -159
rect 453 -160 454 -159
rect 454 -160 455 -159
rect 455 -160 456 -159
rect 456 -160 457 -159
rect 457 -160 458 -159
rect 458 -160 459 -159
rect 459 -160 460 -159
rect 460 -160 461 -159
rect 461 -160 462 -159
rect 462 -160 463 -159
rect 463 -160 464 -159
rect 464 -160 465 -159
rect 465 -160 466 -159
rect 466 -160 467 -159
rect 467 -160 468 -159
rect 468 -160 469 -159
rect 469 -160 470 -159
rect 470 -160 471 -159
rect 471 -160 472 -159
rect 472 -160 473 -159
rect 473 -160 474 -159
rect 474 -160 475 -159
rect 475 -160 476 -159
rect 476 -160 477 -159
rect 477 -160 478 -159
rect 478 -160 479 -159
rect 479 -160 480 -159
rect 2 -161 3 -160
rect 3 -161 4 -160
rect 4 -161 5 -160
rect 5 -161 6 -160
rect 6 -161 7 -160
rect 7 -161 8 -160
rect 8 -161 9 -160
rect 9 -161 10 -160
rect 10 -161 11 -160
rect 11 -161 12 -160
rect 12 -161 13 -160
rect 13 -161 14 -160
rect 14 -161 15 -160
rect 15 -161 16 -160
rect 16 -161 17 -160
rect 17 -161 18 -160
rect 18 -161 19 -160
rect 19 -161 20 -160
rect 20 -161 21 -160
rect 21 -161 22 -160
rect 22 -161 23 -160
rect 23 -161 24 -160
rect 24 -161 25 -160
rect 25 -161 26 -160
rect 26 -161 27 -160
rect 27 -161 28 -160
rect 28 -161 29 -160
rect 29 -161 30 -160
rect 30 -161 31 -160
rect 31 -161 32 -160
rect 32 -161 33 -160
rect 33 -161 34 -160
rect 34 -161 35 -160
rect 35 -161 36 -160
rect 36 -161 37 -160
rect 37 -161 38 -160
rect 38 -161 39 -160
rect 39 -161 40 -160
rect 40 -161 41 -160
rect 41 -161 42 -160
rect 42 -161 43 -160
rect 43 -161 44 -160
rect 44 -161 45 -160
rect 45 -161 46 -160
rect 46 -161 47 -160
rect 47 -161 48 -160
rect 48 -161 49 -160
rect 49 -161 50 -160
rect 50 -161 51 -160
rect 51 -161 52 -160
rect 52 -161 53 -160
rect 53 -161 54 -160
rect 54 -161 55 -160
rect 55 -161 56 -160
rect 56 -161 57 -160
rect 57 -161 58 -160
rect 58 -161 59 -160
rect 59 -161 60 -160
rect 60 -161 61 -160
rect 61 -161 62 -160
rect 62 -161 63 -160
rect 63 -161 64 -160
rect 64 -161 65 -160
rect 65 -161 66 -160
rect 66 -161 67 -160
rect 67 -161 68 -160
rect 68 -161 69 -160
rect 69 -161 70 -160
rect 70 -161 71 -160
rect 71 -161 72 -160
rect 72 -161 73 -160
rect 73 -161 74 -160
rect 74 -161 75 -160
rect 75 -161 76 -160
rect 76 -161 77 -160
rect 77 -161 78 -160
rect 78 -161 79 -160
rect 79 -161 80 -160
rect 80 -161 81 -160
rect 81 -161 82 -160
rect 82 -161 83 -160
rect 83 -161 84 -160
rect 84 -161 85 -160
rect 85 -161 86 -160
rect 86 -161 87 -160
rect 87 -161 88 -160
rect 88 -161 89 -160
rect 89 -161 90 -160
rect 90 -161 91 -160
rect 91 -161 92 -160
rect 92 -161 93 -160
rect 93 -161 94 -160
rect 94 -161 95 -160
rect 95 -161 96 -160
rect 96 -161 97 -160
rect 97 -161 98 -160
rect 98 -161 99 -160
rect 99 -161 100 -160
rect 100 -161 101 -160
rect 101 -161 102 -160
rect 102 -161 103 -160
rect 103 -161 104 -160
rect 104 -161 105 -160
rect 105 -161 106 -160
rect 106 -161 107 -160
rect 107 -161 108 -160
rect 108 -161 109 -160
rect 109 -161 110 -160
rect 110 -161 111 -160
rect 111 -161 112 -160
rect 112 -161 113 -160
rect 113 -161 114 -160
rect 114 -161 115 -160
rect 115 -161 116 -160
rect 116 -161 117 -160
rect 117 -161 118 -160
rect 118 -161 119 -160
rect 119 -161 120 -160
rect 120 -161 121 -160
rect 121 -161 122 -160
rect 122 -161 123 -160
rect 123 -161 124 -160
rect 124 -161 125 -160
rect 125 -161 126 -160
rect 126 -161 127 -160
rect 127 -161 128 -160
rect 128 -161 129 -160
rect 129 -161 130 -160
rect 130 -161 131 -160
rect 131 -161 132 -160
rect 132 -161 133 -160
rect 133 -161 134 -160
rect 134 -161 135 -160
rect 135 -161 136 -160
rect 136 -161 137 -160
rect 137 -161 138 -160
rect 138 -161 139 -160
rect 139 -161 140 -160
rect 140 -161 141 -160
rect 141 -161 142 -160
rect 142 -161 143 -160
rect 143 -161 144 -160
rect 144 -161 145 -160
rect 145 -161 146 -160
rect 146 -161 147 -160
rect 147 -161 148 -160
rect 148 -161 149 -160
rect 149 -161 150 -160
rect 150 -161 151 -160
rect 151 -161 152 -160
rect 152 -161 153 -160
rect 153 -161 154 -160
rect 154 -161 155 -160
rect 155 -161 156 -160
rect 156 -161 157 -160
rect 157 -161 158 -160
rect 158 -161 159 -160
rect 159 -161 160 -160
rect 160 -161 161 -160
rect 161 -161 162 -160
rect 162 -161 163 -160
rect 163 -161 164 -160
rect 164 -161 165 -160
rect 165 -161 166 -160
rect 166 -161 167 -160
rect 167 -161 168 -160
rect 168 -161 169 -160
rect 169 -161 170 -160
rect 170 -161 171 -160
rect 171 -161 172 -160
rect 172 -161 173 -160
rect 173 -161 174 -160
rect 174 -161 175 -160
rect 175 -161 176 -160
rect 176 -161 177 -160
rect 177 -161 178 -160
rect 178 -161 179 -160
rect 179 -161 180 -160
rect 180 -161 181 -160
rect 181 -161 182 -160
rect 182 -161 183 -160
rect 183 -161 184 -160
rect 184 -161 185 -160
rect 185 -161 186 -160
rect 186 -161 187 -160
rect 187 -161 188 -160
rect 188 -161 189 -160
rect 189 -161 190 -160
rect 190 -161 191 -160
rect 191 -161 192 -160
rect 192 -161 193 -160
rect 193 -161 194 -160
rect 194 -161 195 -160
rect 195 -161 196 -160
rect 196 -161 197 -160
rect 197 -161 198 -160
rect 198 -161 199 -160
rect 199 -161 200 -160
rect 200 -161 201 -160
rect 201 -161 202 -160
rect 202 -161 203 -160
rect 203 -161 204 -160
rect 204 -161 205 -160
rect 205 -161 206 -160
rect 206 -161 207 -160
rect 207 -161 208 -160
rect 208 -161 209 -160
rect 209 -161 210 -160
rect 210 -161 211 -160
rect 211 -161 212 -160
rect 212 -161 213 -160
rect 213 -161 214 -160
rect 214 -161 215 -160
rect 215 -161 216 -160
rect 216 -161 217 -160
rect 217 -161 218 -160
rect 218 -161 219 -160
rect 219 -161 220 -160
rect 220 -161 221 -160
rect 221 -161 222 -160
rect 222 -161 223 -160
rect 223 -161 224 -160
rect 224 -161 225 -160
rect 225 -161 226 -160
rect 226 -161 227 -160
rect 227 -161 228 -160
rect 228 -161 229 -160
rect 229 -161 230 -160
rect 230 -161 231 -160
rect 231 -161 232 -160
rect 232 -161 233 -160
rect 233 -161 234 -160
rect 234 -161 235 -160
rect 235 -161 236 -160
rect 236 -161 237 -160
rect 237 -161 238 -160
rect 238 -161 239 -160
rect 239 -161 240 -160
rect 240 -161 241 -160
rect 241 -161 242 -160
rect 242 -161 243 -160
rect 243 -161 244 -160
rect 244 -161 245 -160
rect 245 -161 246 -160
rect 246 -161 247 -160
rect 247 -161 248 -160
rect 248 -161 249 -160
rect 249 -161 250 -160
rect 250 -161 251 -160
rect 251 -161 252 -160
rect 252 -161 253 -160
rect 253 -161 254 -160
rect 254 -161 255 -160
rect 255 -161 256 -160
rect 256 -161 257 -160
rect 257 -161 258 -160
rect 258 -161 259 -160
rect 259 -161 260 -160
rect 260 -161 261 -160
rect 261 -161 262 -160
rect 262 -161 263 -160
rect 263 -161 264 -160
rect 264 -161 265 -160
rect 265 -161 266 -160
rect 266 -161 267 -160
rect 267 -161 268 -160
rect 268 -161 269 -160
rect 269 -161 270 -160
rect 270 -161 271 -160
rect 271 -161 272 -160
rect 272 -161 273 -160
rect 273 -161 274 -160
rect 274 -161 275 -160
rect 275 -161 276 -160
rect 276 -161 277 -160
rect 277 -161 278 -160
rect 278 -161 279 -160
rect 279 -161 280 -160
rect 280 -161 281 -160
rect 281 -161 282 -160
rect 282 -161 283 -160
rect 283 -161 284 -160
rect 284 -161 285 -160
rect 285 -161 286 -160
rect 286 -161 287 -160
rect 287 -161 288 -160
rect 288 -161 289 -160
rect 289 -161 290 -160
rect 290 -161 291 -160
rect 291 -161 292 -160
rect 292 -161 293 -160
rect 293 -161 294 -160
rect 294 -161 295 -160
rect 295 -161 296 -160
rect 296 -161 297 -160
rect 297 -161 298 -160
rect 298 -161 299 -160
rect 299 -161 300 -160
rect 300 -161 301 -160
rect 301 -161 302 -160
rect 302 -161 303 -160
rect 303 -161 304 -160
rect 304 -161 305 -160
rect 305 -161 306 -160
rect 306 -161 307 -160
rect 307 -161 308 -160
rect 308 -161 309 -160
rect 309 -161 310 -160
rect 310 -161 311 -160
rect 311 -161 312 -160
rect 312 -161 313 -160
rect 313 -161 314 -160
rect 314 -161 315 -160
rect 315 -161 316 -160
rect 316 -161 317 -160
rect 317 -161 318 -160
rect 318 -161 319 -160
rect 319 -161 320 -160
rect 320 -161 321 -160
rect 321 -161 322 -160
rect 322 -161 323 -160
rect 323 -161 324 -160
rect 324 -161 325 -160
rect 325 -161 326 -160
rect 326 -161 327 -160
rect 327 -161 328 -160
rect 328 -161 329 -160
rect 329 -161 330 -160
rect 330 -161 331 -160
rect 331 -161 332 -160
rect 332 -161 333 -160
rect 333 -161 334 -160
rect 334 -161 335 -160
rect 335 -161 336 -160
rect 336 -161 337 -160
rect 337 -161 338 -160
rect 338 -161 339 -160
rect 339 -161 340 -160
rect 340 -161 341 -160
rect 341 -161 342 -160
rect 342 -161 343 -160
rect 343 -161 344 -160
rect 344 -161 345 -160
rect 345 -161 346 -160
rect 346 -161 347 -160
rect 347 -161 348 -160
rect 348 -161 349 -160
rect 349 -161 350 -160
rect 350 -161 351 -160
rect 351 -161 352 -160
rect 352 -161 353 -160
rect 353 -161 354 -160
rect 354 -161 355 -160
rect 355 -161 356 -160
rect 356 -161 357 -160
rect 357 -161 358 -160
rect 358 -161 359 -160
rect 359 -161 360 -160
rect 360 -161 361 -160
rect 361 -161 362 -160
rect 362 -161 363 -160
rect 363 -161 364 -160
rect 364 -161 365 -160
rect 365 -161 366 -160
rect 366 -161 367 -160
rect 367 -161 368 -160
rect 368 -161 369 -160
rect 369 -161 370 -160
rect 370 -161 371 -160
rect 371 -161 372 -160
rect 372 -161 373 -160
rect 373 -161 374 -160
rect 374 -161 375 -160
rect 375 -161 376 -160
rect 376 -161 377 -160
rect 377 -161 378 -160
rect 378 -161 379 -160
rect 379 -161 380 -160
rect 380 -161 381 -160
rect 381 -161 382 -160
rect 382 -161 383 -160
rect 383 -161 384 -160
rect 384 -161 385 -160
rect 385 -161 386 -160
rect 386 -161 387 -160
rect 387 -161 388 -160
rect 388 -161 389 -160
rect 389 -161 390 -160
rect 390 -161 391 -160
rect 391 -161 392 -160
rect 392 -161 393 -160
rect 393 -161 394 -160
rect 394 -161 395 -160
rect 395 -161 396 -160
rect 396 -161 397 -160
rect 397 -161 398 -160
rect 398 -161 399 -160
rect 399 -161 400 -160
rect 400 -161 401 -160
rect 401 -161 402 -160
rect 402 -161 403 -160
rect 403 -161 404 -160
rect 404 -161 405 -160
rect 405 -161 406 -160
rect 406 -161 407 -160
rect 407 -161 408 -160
rect 408 -161 409 -160
rect 409 -161 410 -160
rect 410 -161 411 -160
rect 411 -161 412 -160
rect 412 -161 413 -160
rect 413 -161 414 -160
rect 414 -161 415 -160
rect 415 -161 416 -160
rect 416 -161 417 -160
rect 417 -161 418 -160
rect 418 -161 419 -160
rect 419 -161 420 -160
rect 420 -161 421 -160
rect 421 -161 422 -160
rect 422 -161 423 -160
rect 423 -161 424 -160
rect 424 -161 425 -160
rect 425 -161 426 -160
rect 426 -161 427 -160
rect 427 -161 428 -160
rect 428 -161 429 -160
rect 429 -161 430 -160
rect 430 -161 431 -160
rect 431 -161 432 -160
rect 432 -161 433 -160
rect 433 -161 434 -160
rect 434 -161 435 -160
rect 435 -161 436 -160
rect 436 -161 437 -160
rect 437 -161 438 -160
rect 438 -161 439 -160
rect 439 -161 440 -160
rect 440 -161 441 -160
rect 441 -161 442 -160
rect 442 -161 443 -160
rect 443 -161 444 -160
rect 444 -161 445 -160
rect 445 -161 446 -160
rect 446 -161 447 -160
rect 447 -161 448 -160
rect 448 -161 449 -160
rect 449 -161 450 -160
rect 450 -161 451 -160
rect 451 -161 452 -160
rect 452 -161 453 -160
rect 453 -161 454 -160
rect 454 -161 455 -160
rect 455 -161 456 -160
rect 456 -161 457 -160
rect 457 -161 458 -160
rect 458 -161 459 -160
rect 459 -161 460 -160
rect 460 -161 461 -160
rect 461 -161 462 -160
rect 462 -161 463 -160
rect 463 -161 464 -160
rect 464 -161 465 -160
rect 465 -161 466 -160
rect 466 -161 467 -160
rect 467 -161 468 -160
rect 468 -161 469 -160
rect 469 -161 470 -160
rect 470 -161 471 -160
rect 471 -161 472 -160
rect 472 -161 473 -160
rect 473 -161 474 -160
rect 474 -161 475 -160
rect 475 -161 476 -160
rect 476 -161 477 -160
rect 477 -161 478 -160
rect 478 -161 479 -160
rect 479 -161 480 -160
rect 2 -162 3 -161
rect 3 -162 4 -161
rect 4 -162 5 -161
rect 5 -162 6 -161
rect 6 -162 7 -161
rect 7 -162 8 -161
rect 8 -162 9 -161
rect 9 -162 10 -161
rect 10 -162 11 -161
rect 11 -162 12 -161
rect 12 -162 13 -161
rect 13 -162 14 -161
rect 14 -162 15 -161
rect 15 -162 16 -161
rect 16 -162 17 -161
rect 17 -162 18 -161
rect 18 -162 19 -161
rect 19 -162 20 -161
rect 20 -162 21 -161
rect 21 -162 22 -161
rect 22 -162 23 -161
rect 23 -162 24 -161
rect 24 -162 25 -161
rect 25 -162 26 -161
rect 26 -162 27 -161
rect 27 -162 28 -161
rect 28 -162 29 -161
rect 29 -162 30 -161
rect 30 -162 31 -161
rect 31 -162 32 -161
rect 32 -162 33 -161
rect 33 -162 34 -161
rect 34 -162 35 -161
rect 35 -162 36 -161
rect 36 -162 37 -161
rect 37 -162 38 -161
rect 38 -162 39 -161
rect 39 -162 40 -161
rect 40 -162 41 -161
rect 41 -162 42 -161
rect 42 -162 43 -161
rect 43 -162 44 -161
rect 44 -162 45 -161
rect 45 -162 46 -161
rect 46 -162 47 -161
rect 47 -162 48 -161
rect 48 -162 49 -161
rect 49 -162 50 -161
rect 50 -162 51 -161
rect 51 -162 52 -161
rect 52 -162 53 -161
rect 53 -162 54 -161
rect 54 -162 55 -161
rect 55 -162 56 -161
rect 56 -162 57 -161
rect 57 -162 58 -161
rect 58 -162 59 -161
rect 59 -162 60 -161
rect 60 -162 61 -161
rect 61 -162 62 -161
rect 62 -162 63 -161
rect 63 -162 64 -161
rect 64 -162 65 -161
rect 65 -162 66 -161
rect 66 -162 67 -161
rect 67 -162 68 -161
rect 68 -162 69 -161
rect 69 -162 70 -161
rect 70 -162 71 -161
rect 71 -162 72 -161
rect 72 -162 73 -161
rect 73 -162 74 -161
rect 74 -162 75 -161
rect 75 -162 76 -161
rect 76 -162 77 -161
rect 77 -162 78 -161
rect 78 -162 79 -161
rect 79 -162 80 -161
rect 80 -162 81 -161
rect 81 -162 82 -161
rect 82 -162 83 -161
rect 83 -162 84 -161
rect 84 -162 85 -161
rect 85 -162 86 -161
rect 86 -162 87 -161
rect 87 -162 88 -161
rect 88 -162 89 -161
rect 89 -162 90 -161
rect 90 -162 91 -161
rect 91 -162 92 -161
rect 92 -162 93 -161
rect 93 -162 94 -161
rect 94 -162 95 -161
rect 95 -162 96 -161
rect 96 -162 97 -161
rect 97 -162 98 -161
rect 98 -162 99 -161
rect 99 -162 100 -161
rect 100 -162 101 -161
rect 101 -162 102 -161
rect 102 -162 103 -161
rect 103 -162 104 -161
rect 104 -162 105 -161
rect 105 -162 106 -161
rect 106 -162 107 -161
rect 107 -162 108 -161
rect 108 -162 109 -161
rect 109 -162 110 -161
rect 110 -162 111 -161
rect 111 -162 112 -161
rect 112 -162 113 -161
rect 113 -162 114 -161
rect 114 -162 115 -161
rect 115 -162 116 -161
rect 116 -162 117 -161
rect 117 -162 118 -161
rect 118 -162 119 -161
rect 119 -162 120 -161
rect 120 -162 121 -161
rect 121 -162 122 -161
rect 122 -162 123 -161
rect 123 -162 124 -161
rect 124 -162 125 -161
rect 125 -162 126 -161
rect 126 -162 127 -161
rect 127 -162 128 -161
rect 128 -162 129 -161
rect 129 -162 130 -161
rect 130 -162 131 -161
rect 131 -162 132 -161
rect 132 -162 133 -161
rect 133 -162 134 -161
rect 134 -162 135 -161
rect 135 -162 136 -161
rect 136 -162 137 -161
rect 137 -162 138 -161
rect 138 -162 139 -161
rect 139 -162 140 -161
rect 140 -162 141 -161
rect 141 -162 142 -161
rect 142 -162 143 -161
rect 143 -162 144 -161
rect 144 -162 145 -161
rect 145 -162 146 -161
rect 146 -162 147 -161
rect 147 -162 148 -161
rect 148 -162 149 -161
rect 149 -162 150 -161
rect 150 -162 151 -161
rect 151 -162 152 -161
rect 152 -162 153 -161
rect 153 -162 154 -161
rect 154 -162 155 -161
rect 155 -162 156 -161
rect 156 -162 157 -161
rect 157 -162 158 -161
rect 158 -162 159 -161
rect 159 -162 160 -161
rect 160 -162 161 -161
rect 161 -162 162 -161
rect 162 -162 163 -161
rect 163 -162 164 -161
rect 164 -162 165 -161
rect 165 -162 166 -161
rect 166 -162 167 -161
rect 167 -162 168 -161
rect 168 -162 169 -161
rect 169 -162 170 -161
rect 170 -162 171 -161
rect 171 -162 172 -161
rect 172 -162 173 -161
rect 173 -162 174 -161
rect 174 -162 175 -161
rect 175 -162 176 -161
rect 176 -162 177 -161
rect 177 -162 178 -161
rect 178 -162 179 -161
rect 179 -162 180 -161
rect 180 -162 181 -161
rect 181 -162 182 -161
rect 182 -162 183 -161
rect 183 -162 184 -161
rect 184 -162 185 -161
rect 185 -162 186 -161
rect 186 -162 187 -161
rect 187 -162 188 -161
rect 188 -162 189 -161
rect 189 -162 190 -161
rect 190 -162 191 -161
rect 191 -162 192 -161
rect 192 -162 193 -161
rect 193 -162 194 -161
rect 194 -162 195 -161
rect 195 -162 196 -161
rect 196 -162 197 -161
rect 197 -162 198 -161
rect 198 -162 199 -161
rect 199 -162 200 -161
rect 200 -162 201 -161
rect 201 -162 202 -161
rect 202 -162 203 -161
rect 203 -162 204 -161
rect 204 -162 205 -161
rect 205 -162 206 -161
rect 206 -162 207 -161
rect 207 -162 208 -161
rect 208 -162 209 -161
rect 209 -162 210 -161
rect 210 -162 211 -161
rect 211 -162 212 -161
rect 212 -162 213 -161
rect 213 -162 214 -161
rect 214 -162 215 -161
rect 215 -162 216 -161
rect 216 -162 217 -161
rect 217 -162 218 -161
rect 218 -162 219 -161
rect 219 -162 220 -161
rect 220 -162 221 -161
rect 221 -162 222 -161
rect 222 -162 223 -161
rect 223 -162 224 -161
rect 224 -162 225 -161
rect 225 -162 226 -161
rect 226 -162 227 -161
rect 227 -162 228 -161
rect 228 -162 229 -161
rect 229 -162 230 -161
rect 230 -162 231 -161
rect 231 -162 232 -161
rect 232 -162 233 -161
rect 233 -162 234 -161
rect 234 -162 235 -161
rect 235 -162 236 -161
rect 236 -162 237 -161
rect 237 -162 238 -161
rect 238 -162 239 -161
rect 239 -162 240 -161
rect 240 -162 241 -161
rect 241 -162 242 -161
rect 242 -162 243 -161
rect 243 -162 244 -161
rect 244 -162 245 -161
rect 245 -162 246 -161
rect 246 -162 247 -161
rect 247 -162 248 -161
rect 248 -162 249 -161
rect 249 -162 250 -161
rect 250 -162 251 -161
rect 251 -162 252 -161
rect 252 -162 253 -161
rect 253 -162 254 -161
rect 254 -162 255 -161
rect 255 -162 256 -161
rect 256 -162 257 -161
rect 257 -162 258 -161
rect 258 -162 259 -161
rect 259 -162 260 -161
rect 260 -162 261 -161
rect 261 -162 262 -161
rect 262 -162 263 -161
rect 263 -162 264 -161
rect 264 -162 265 -161
rect 265 -162 266 -161
rect 266 -162 267 -161
rect 267 -162 268 -161
rect 268 -162 269 -161
rect 269 -162 270 -161
rect 270 -162 271 -161
rect 271 -162 272 -161
rect 272 -162 273 -161
rect 273 -162 274 -161
rect 274 -162 275 -161
rect 275 -162 276 -161
rect 276 -162 277 -161
rect 277 -162 278 -161
rect 278 -162 279 -161
rect 279 -162 280 -161
rect 280 -162 281 -161
rect 281 -162 282 -161
rect 282 -162 283 -161
rect 283 -162 284 -161
rect 284 -162 285 -161
rect 285 -162 286 -161
rect 286 -162 287 -161
rect 287 -162 288 -161
rect 288 -162 289 -161
rect 289 -162 290 -161
rect 290 -162 291 -161
rect 291 -162 292 -161
rect 292 -162 293 -161
rect 293 -162 294 -161
rect 294 -162 295 -161
rect 295 -162 296 -161
rect 296 -162 297 -161
rect 297 -162 298 -161
rect 298 -162 299 -161
rect 299 -162 300 -161
rect 300 -162 301 -161
rect 301 -162 302 -161
rect 302 -162 303 -161
rect 303 -162 304 -161
rect 304 -162 305 -161
rect 305 -162 306 -161
rect 306 -162 307 -161
rect 307 -162 308 -161
rect 308 -162 309 -161
rect 309 -162 310 -161
rect 310 -162 311 -161
rect 311 -162 312 -161
rect 312 -162 313 -161
rect 313 -162 314 -161
rect 314 -162 315 -161
rect 315 -162 316 -161
rect 316 -162 317 -161
rect 317 -162 318 -161
rect 318 -162 319 -161
rect 319 -162 320 -161
rect 320 -162 321 -161
rect 321 -162 322 -161
rect 322 -162 323 -161
rect 323 -162 324 -161
rect 324 -162 325 -161
rect 325 -162 326 -161
rect 326 -162 327 -161
rect 327 -162 328 -161
rect 328 -162 329 -161
rect 329 -162 330 -161
rect 330 -162 331 -161
rect 331 -162 332 -161
rect 332 -162 333 -161
rect 333 -162 334 -161
rect 334 -162 335 -161
rect 335 -162 336 -161
rect 336 -162 337 -161
rect 337 -162 338 -161
rect 338 -162 339 -161
rect 339 -162 340 -161
rect 340 -162 341 -161
rect 341 -162 342 -161
rect 342 -162 343 -161
rect 343 -162 344 -161
rect 344 -162 345 -161
rect 345 -162 346 -161
rect 346 -162 347 -161
rect 347 -162 348 -161
rect 348 -162 349 -161
rect 349 -162 350 -161
rect 350 -162 351 -161
rect 351 -162 352 -161
rect 352 -162 353 -161
rect 353 -162 354 -161
rect 354 -162 355 -161
rect 355 -162 356 -161
rect 356 -162 357 -161
rect 357 -162 358 -161
rect 358 -162 359 -161
rect 359 -162 360 -161
rect 360 -162 361 -161
rect 361 -162 362 -161
rect 362 -162 363 -161
rect 363 -162 364 -161
rect 364 -162 365 -161
rect 365 -162 366 -161
rect 366 -162 367 -161
rect 367 -162 368 -161
rect 368 -162 369 -161
rect 369 -162 370 -161
rect 370 -162 371 -161
rect 371 -162 372 -161
rect 372 -162 373 -161
rect 373 -162 374 -161
rect 374 -162 375 -161
rect 375 -162 376 -161
rect 376 -162 377 -161
rect 377 -162 378 -161
rect 378 -162 379 -161
rect 379 -162 380 -161
rect 380 -162 381 -161
rect 381 -162 382 -161
rect 382 -162 383 -161
rect 383 -162 384 -161
rect 384 -162 385 -161
rect 385 -162 386 -161
rect 386 -162 387 -161
rect 387 -162 388 -161
rect 388 -162 389 -161
rect 389 -162 390 -161
rect 390 -162 391 -161
rect 391 -162 392 -161
rect 392 -162 393 -161
rect 393 -162 394 -161
rect 394 -162 395 -161
rect 395 -162 396 -161
rect 396 -162 397 -161
rect 397 -162 398 -161
rect 398 -162 399 -161
rect 399 -162 400 -161
rect 400 -162 401 -161
rect 401 -162 402 -161
rect 402 -162 403 -161
rect 403 -162 404 -161
rect 404 -162 405 -161
rect 405 -162 406 -161
rect 406 -162 407 -161
rect 407 -162 408 -161
rect 408 -162 409 -161
rect 409 -162 410 -161
rect 410 -162 411 -161
rect 411 -162 412 -161
rect 412 -162 413 -161
rect 413 -162 414 -161
rect 414 -162 415 -161
rect 415 -162 416 -161
rect 416 -162 417 -161
rect 417 -162 418 -161
rect 418 -162 419 -161
rect 419 -162 420 -161
rect 420 -162 421 -161
rect 421 -162 422 -161
rect 422 -162 423 -161
rect 423 -162 424 -161
rect 424 -162 425 -161
rect 425 -162 426 -161
rect 426 -162 427 -161
rect 427 -162 428 -161
rect 428 -162 429 -161
rect 429 -162 430 -161
rect 430 -162 431 -161
rect 431 -162 432 -161
rect 432 -162 433 -161
rect 433 -162 434 -161
rect 434 -162 435 -161
rect 435 -162 436 -161
rect 436 -162 437 -161
rect 437 -162 438 -161
rect 438 -162 439 -161
rect 439 -162 440 -161
rect 440 -162 441 -161
rect 441 -162 442 -161
rect 442 -162 443 -161
rect 443 -162 444 -161
rect 444 -162 445 -161
rect 445 -162 446 -161
rect 446 -162 447 -161
rect 447 -162 448 -161
rect 448 -162 449 -161
rect 449 -162 450 -161
rect 450 -162 451 -161
rect 451 -162 452 -161
rect 452 -162 453 -161
rect 453 -162 454 -161
rect 454 -162 455 -161
rect 455 -162 456 -161
rect 456 -162 457 -161
rect 457 -162 458 -161
rect 458 -162 459 -161
rect 459 -162 460 -161
rect 460 -162 461 -161
rect 461 -162 462 -161
rect 462 -162 463 -161
rect 463 -162 464 -161
rect 464 -162 465 -161
rect 465 -162 466 -161
rect 466 -162 467 -161
rect 467 -162 468 -161
rect 468 -162 469 -161
rect 469 -162 470 -161
rect 470 -162 471 -161
rect 471 -162 472 -161
rect 472 -162 473 -161
rect 473 -162 474 -161
rect 474 -162 475 -161
rect 475 -162 476 -161
rect 476 -162 477 -161
rect 477 -162 478 -161
rect 478 -162 479 -161
rect 479 -162 480 -161
rect 2 -163 3 -162
rect 3 -163 4 -162
rect 4 -163 5 -162
rect 5 -163 6 -162
rect 6 -163 7 -162
rect 7 -163 8 -162
rect 8 -163 9 -162
rect 9 -163 10 -162
rect 10 -163 11 -162
rect 11 -163 12 -162
rect 12 -163 13 -162
rect 13 -163 14 -162
rect 14 -163 15 -162
rect 15 -163 16 -162
rect 16 -163 17 -162
rect 17 -163 18 -162
rect 18 -163 19 -162
rect 19 -163 20 -162
rect 20 -163 21 -162
rect 21 -163 22 -162
rect 22 -163 23 -162
rect 23 -163 24 -162
rect 24 -163 25 -162
rect 25 -163 26 -162
rect 26 -163 27 -162
rect 27 -163 28 -162
rect 28 -163 29 -162
rect 29 -163 30 -162
rect 30 -163 31 -162
rect 31 -163 32 -162
rect 32 -163 33 -162
rect 33 -163 34 -162
rect 34 -163 35 -162
rect 35 -163 36 -162
rect 36 -163 37 -162
rect 37 -163 38 -162
rect 38 -163 39 -162
rect 39 -163 40 -162
rect 40 -163 41 -162
rect 41 -163 42 -162
rect 42 -163 43 -162
rect 43 -163 44 -162
rect 44 -163 45 -162
rect 45 -163 46 -162
rect 46 -163 47 -162
rect 47 -163 48 -162
rect 48 -163 49 -162
rect 49 -163 50 -162
rect 50 -163 51 -162
rect 51 -163 52 -162
rect 52 -163 53 -162
rect 53 -163 54 -162
rect 54 -163 55 -162
rect 55 -163 56 -162
rect 56 -163 57 -162
rect 57 -163 58 -162
rect 58 -163 59 -162
rect 59 -163 60 -162
rect 60 -163 61 -162
rect 61 -163 62 -162
rect 62 -163 63 -162
rect 63 -163 64 -162
rect 64 -163 65 -162
rect 65 -163 66 -162
rect 66 -163 67 -162
rect 67 -163 68 -162
rect 68 -163 69 -162
rect 69 -163 70 -162
rect 70 -163 71 -162
rect 71 -163 72 -162
rect 72 -163 73 -162
rect 73 -163 74 -162
rect 74 -163 75 -162
rect 75 -163 76 -162
rect 76 -163 77 -162
rect 77 -163 78 -162
rect 78 -163 79 -162
rect 79 -163 80 -162
rect 80 -163 81 -162
rect 81 -163 82 -162
rect 82 -163 83 -162
rect 83 -163 84 -162
rect 84 -163 85 -162
rect 85 -163 86 -162
rect 86 -163 87 -162
rect 87 -163 88 -162
rect 88 -163 89 -162
rect 89 -163 90 -162
rect 90 -163 91 -162
rect 91 -163 92 -162
rect 92 -163 93 -162
rect 93 -163 94 -162
rect 94 -163 95 -162
rect 95 -163 96 -162
rect 96 -163 97 -162
rect 97 -163 98 -162
rect 98 -163 99 -162
rect 99 -163 100 -162
rect 100 -163 101 -162
rect 101 -163 102 -162
rect 102 -163 103 -162
rect 103 -163 104 -162
rect 104 -163 105 -162
rect 105 -163 106 -162
rect 106 -163 107 -162
rect 107 -163 108 -162
rect 108 -163 109 -162
rect 109 -163 110 -162
rect 110 -163 111 -162
rect 111 -163 112 -162
rect 112 -163 113 -162
rect 113 -163 114 -162
rect 114 -163 115 -162
rect 115 -163 116 -162
rect 116 -163 117 -162
rect 117 -163 118 -162
rect 118 -163 119 -162
rect 119 -163 120 -162
rect 120 -163 121 -162
rect 121 -163 122 -162
rect 122 -163 123 -162
rect 123 -163 124 -162
rect 124 -163 125 -162
rect 125 -163 126 -162
rect 126 -163 127 -162
rect 127 -163 128 -162
rect 128 -163 129 -162
rect 129 -163 130 -162
rect 130 -163 131 -162
rect 131 -163 132 -162
rect 132 -163 133 -162
rect 133 -163 134 -162
rect 134 -163 135 -162
rect 135 -163 136 -162
rect 136 -163 137 -162
rect 137 -163 138 -162
rect 138 -163 139 -162
rect 139 -163 140 -162
rect 140 -163 141 -162
rect 141 -163 142 -162
rect 142 -163 143 -162
rect 143 -163 144 -162
rect 144 -163 145 -162
rect 145 -163 146 -162
rect 146 -163 147 -162
rect 147 -163 148 -162
rect 148 -163 149 -162
rect 149 -163 150 -162
rect 150 -163 151 -162
rect 151 -163 152 -162
rect 152 -163 153 -162
rect 153 -163 154 -162
rect 154 -163 155 -162
rect 155 -163 156 -162
rect 156 -163 157 -162
rect 157 -163 158 -162
rect 158 -163 159 -162
rect 159 -163 160 -162
rect 160 -163 161 -162
rect 161 -163 162 -162
rect 162 -163 163 -162
rect 163 -163 164 -162
rect 164 -163 165 -162
rect 165 -163 166 -162
rect 166 -163 167 -162
rect 167 -163 168 -162
rect 168 -163 169 -162
rect 169 -163 170 -162
rect 170 -163 171 -162
rect 171 -163 172 -162
rect 172 -163 173 -162
rect 173 -163 174 -162
rect 174 -163 175 -162
rect 175 -163 176 -162
rect 176 -163 177 -162
rect 177 -163 178 -162
rect 178 -163 179 -162
rect 179 -163 180 -162
rect 180 -163 181 -162
rect 181 -163 182 -162
rect 182 -163 183 -162
rect 183 -163 184 -162
rect 184 -163 185 -162
rect 185 -163 186 -162
rect 186 -163 187 -162
rect 187 -163 188 -162
rect 188 -163 189 -162
rect 189 -163 190 -162
rect 190 -163 191 -162
rect 191 -163 192 -162
rect 192 -163 193 -162
rect 193 -163 194 -162
rect 194 -163 195 -162
rect 195 -163 196 -162
rect 196 -163 197 -162
rect 197 -163 198 -162
rect 198 -163 199 -162
rect 199 -163 200 -162
rect 200 -163 201 -162
rect 201 -163 202 -162
rect 202 -163 203 -162
rect 203 -163 204 -162
rect 204 -163 205 -162
rect 205 -163 206 -162
rect 206 -163 207 -162
rect 207 -163 208 -162
rect 208 -163 209 -162
rect 209 -163 210 -162
rect 210 -163 211 -162
rect 211 -163 212 -162
rect 212 -163 213 -162
rect 213 -163 214 -162
rect 214 -163 215 -162
rect 215 -163 216 -162
rect 216 -163 217 -162
rect 217 -163 218 -162
rect 218 -163 219 -162
rect 219 -163 220 -162
rect 220 -163 221 -162
rect 221 -163 222 -162
rect 222 -163 223 -162
rect 223 -163 224 -162
rect 224 -163 225 -162
rect 225 -163 226 -162
rect 226 -163 227 -162
rect 227 -163 228 -162
rect 228 -163 229 -162
rect 229 -163 230 -162
rect 230 -163 231 -162
rect 231 -163 232 -162
rect 232 -163 233 -162
rect 233 -163 234 -162
rect 234 -163 235 -162
rect 235 -163 236 -162
rect 236 -163 237 -162
rect 237 -163 238 -162
rect 238 -163 239 -162
rect 239 -163 240 -162
rect 240 -163 241 -162
rect 241 -163 242 -162
rect 242 -163 243 -162
rect 243 -163 244 -162
rect 244 -163 245 -162
rect 245 -163 246 -162
rect 246 -163 247 -162
rect 247 -163 248 -162
rect 248 -163 249 -162
rect 249 -163 250 -162
rect 250 -163 251 -162
rect 251 -163 252 -162
rect 252 -163 253 -162
rect 253 -163 254 -162
rect 254 -163 255 -162
rect 255 -163 256 -162
rect 256 -163 257 -162
rect 257 -163 258 -162
rect 258 -163 259 -162
rect 259 -163 260 -162
rect 260 -163 261 -162
rect 261 -163 262 -162
rect 262 -163 263 -162
rect 263 -163 264 -162
rect 264 -163 265 -162
rect 265 -163 266 -162
rect 266 -163 267 -162
rect 267 -163 268 -162
rect 268 -163 269 -162
rect 269 -163 270 -162
rect 270 -163 271 -162
rect 271 -163 272 -162
rect 272 -163 273 -162
rect 273 -163 274 -162
rect 274 -163 275 -162
rect 275 -163 276 -162
rect 276 -163 277 -162
rect 277 -163 278 -162
rect 278 -163 279 -162
rect 279 -163 280 -162
rect 280 -163 281 -162
rect 281 -163 282 -162
rect 282 -163 283 -162
rect 283 -163 284 -162
rect 284 -163 285 -162
rect 285 -163 286 -162
rect 286 -163 287 -162
rect 287 -163 288 -162
rect 288 -163 289 -162
rect 289 -163 290 -162
rect 290 -163 291 -162
rect 291 -163 292 -162
rect 292 -163 293 -162
rect 293 -163 294 -162
rect 294 -163 295 -162
rect 295 -163 296 -162
rect 296 -163 297 -162
rect 297 -163 298 -162
rect 298 -163 299 -162
rect 299 -163 300 -162
rect 300 -163 301 -162
rect 301 -163 302 -162
rect 302 -163 303 -162
rect 303 -163 304 -162
rect 304 -163 305 -162
rect 305 -163 306 -162
rect 306 -163 307 -162
rect 307 -163 308 -162
rect 308 -163 309 -162
rect 309 -163 310 -162
rect 310 -163 311 -162
rect 311 -163 312 -162
rect 312 -163 313 -162
rect 313 -163 314 -162
rect 314 -163 315 -162
rect 315 -163 316 -162
rect 316 -163 317 -162
rect 317 -163 318 -162
rect 318 -163 319 -162
rect 319 -163 320 -162
rect 320 -163 321 -162
rect 321 -163 322 -162
rect 322 -163 323 -162
rect 323 -163 324 -162
rect 324 -163 325 -162
rect 325 -163 326 -162
rect 326 -163 327 -162
rect 327 -163 328 -162
rect 328 -163 329 -162
rect 329 -163 330 -162
rect 330 -163 331 -162
rect 331 -163 332 -162
rect 332 -163 333 -162
rect 333 -163 334 -162
rect 334 -163 335 -162
rect 335 -163 336 -162
rect 336 -163 337 -162
rect 337 -163 338 -162
rect 338 -163 339 -162
rect 339 -163 340 -162
rect 340 -163 341 -162
rect 341 -163 342 -162
rect 342 -163 343 -162
rect 343 -163 344 -162
rect 344 -163 345 -162
rect 345 -163 346 -162
rect 346 -163 347 -162
rect 347 -163 348 -162
rect 348 -163 349 -162
rect 349 -163 350 -162
rect 350 -163 351 -162
rect 351 -163 352 -162
rect 352 -163 353 -162
rect 353 -163 354 -162
rect 354 -163 355 -162
rect 355 -163 356 -162
rect 356 -163 357 -162
rect 357 -163 358 -162
rect 358 -163 359 -162
rect 359 -163 360 -162
rect 360 -163 361 -162
rect 361 -163 362 -162
rect 362 -163 363 -162
rect 363 -163 364 -162
rect 364 -163 365 -162
rect 365 -163 366 -162
rect 366 -163 367 -162
rect 367 -163 368 -162
rect 368 -163 369 -162
rect 369 -163 370 -162
rect 370 -163 371 -162
rect 371 -163 372 -162
rect 372 -163 373 -162
rect 373 -163 374 -162
rect 374 -163 375 -162
rect 375 -163 376 -162
rect 376 -163 377 -162
rect 377 -163 378 -162
rect 378 -163 379 -162
rect 379 -163 380 -162
rect 380 -163 381 -162
rect 381 -163 382 -162
rect 382 -163 383 -162
rect 383 -163 384 -162
rect 384 -163 385 -162
rect 385 -163 386 -162
rect 386 -163 387 -162
rect 387 -163 388 -162
rect 388 -163 389 -162
rect 389 -163 390 -162
rect 390 -163 391 -162
rect 391 -163 392 -162
rect 392 -163 393 -162
rect 393 -163 394 -162
rect 394 -163 395 -162
rect 395 -163 396 -162
rect 396 -163 397 -162
rect 397 -163 398 -162
rect 398 -163 399 -162
rect 399 -163 400 -162
rect 400 -163 401 -162
rect 401 -163 402 -162
rect 402 -163 403 -162
rect 403 -163 404 -162
rect 404 -163 405 -162
rect 405 -163 406 -162
rect 406 -163 407 -162
rect 407 -163 408 -162
rect 408 -163 409 -162
rect 409 -163 410 -162
rect 410 -163 411 -162
rect 411 -163 412 -162
rect 412 -163 413 -162
rect 413 -163 414 -162
rect 414 -163 415 -162
rect 415 -163 416 -162
rect 416 -163 417 -162
rect 417 -163 418 -162
rect 418 -163 419 -162
rect 419 -163 420 -162
rect 420 -163 421 -162
rect 421 -163 422 -162
rect 422 -163 423 -162
rect 423 -163 424 -162
rect 424 -163 425 -162
rect 425 -163 426 -162
rect 426 -163 427 -162
rect 427 -163 428 -162
rect 428 -163 429 -162
rect 429 -163 430 -162
rect 430 -163 431 -162
rect 431 -163 432 -162
rect 432 -163 433 -162
rect 433 -163 434 -162
rect 434 -163 435 -162
rect 435 -163 436 -162
rect 436 -163 437 -162
rect 437 -163 438 -162
rect 438 -163 439 -162
rect 439 -163 440 -162
rect 440 -163 441 -162
rect 441 -163 442 -162
rect 442 -163 443 -162
rect 443 -163 444 -162
rect 444 -163 445 -162
rect 445 -163 446 -162
rect 446 -163 447 -162
rect 447 -163 448 -162
rect 448 -163 449 -162
rect 449 -163 450 -162
rect 450 -163 451 -162
rect 451 -163 452 -162
rect 452 -163 453 -162
rect 453 -163 454 -162
rect 454 -163 455 -162
rect 455 -163 456 -162
rect 456 -163 457 -162
rect 457 -163 458 -162
rect 458 -163 459 -162
rect 459 -163 460 -162
rect 460 -163 461 -162
rect 461 -163 462 -162
rect 462 -163 463 -162
rect 463 -163 464 -162
rect 464 -163 465 -162
rect 465 -163 466 -162
rect 466 -163 467 -162
rect 467 -163 468 -162
rect 468 -163 469 -162
rect 469 -163 470 -162
rect 470 -163 471 -162
rect 471 -163 472 -162
rect 472 -163 473 -162
rect 473 -163 474 -162
rect 474 -163 475 -162
rect 475 -163 476 -162
rect 476 -163 477 -162
rect 477 -163 478 -162
rect 478 -163 479 -162
rect 479 -163 480 -162
rect 2 -164 3 -163
rect 3 -164 4 -163
rect 4 -164 5 -163
rect 5 -164 6 -163
rect 6 -164 7 -163
rect 7 -164 8 -163
rect 8 -164 9 -163
rect 9 -164 10 -163
rect 10 -164 11 -163
rect 11 -164 12 -163
rect 12 -164 13 -163
rect 13 -164 14 -163
rect 14 -164 15 -163
rect 15 -164 16 -163
rect 16 -164 17 -163
rect 17 -164 18 -163
rect 18 -164 19 -163
rect 19 -164 20 -163
rect 20 -164 21 -163
rect 21 -164 22 -163
rect 22 -164 23 -163
rect 23 -164 24 -163
rect 24 -164 25 -163
rect 25 -164 26 -163
rect 26 -164 27 -163
rect 27 -164 28 -163
rect 28 -164 29 -163
rect 29 -164 30 -163
rect 30 -164 31 -163
rect 31 -164 32 -163
rect 32 -164 33 -163
rect 33 -164 34 -163
rect 34 -164 35 -163
rect 35 -164 36 -163
rect 36 -164 37 -163
rect 37 -164 38 -163
rect 38 -164 39 -163
rect 39 -164 40 -163
rect 40 -164 41 -163
rect 41 -164 42 -163
rect 42 -164 43 -163
rect 43 -164 44 -163
rect 44 -164 45 -163
rect 45 -164 46 -163
rect 46 -164 47 -163
rect 47 -164 48 -163
rect 48 -164 49 -163
rect 49 -164 50 -163
rect 50 -164 51 -163
rect 51 -164 52 -163
rect 52 -164 53 -163
rect 53 -164 54 -163
rect 54 -164 55 -163
rect 55 -164 56 -163
rect 56 -164 57 -163
rect 57 -164 58 -163
rect 58 -164 59 -163
rect 59 -164 60 -163
rect 60 -164 61 -163
rect 61 -164 62 -163
rect 62 -164 63 -163
rect 63 -164 64 -163
rect 64 -164 65 -163
rect 65 -164 66 -163
rect 66 -164 67 -163
rect 67 -164 68 -163
rect 68 -164 69 -163
rect 69 -164 70 -163
rect 70 -164 71 -163
rect 71 -164 72 -163
rect 72 -164 73 -163
rect 73 -164 74 -163
rect 74 -164 75 -163
rect 75 -164 76 -163
rect 76 -164 77 -163
rect 77 -164 78 -163
rect 78 -164 79 -163
rect 79 -164 80 -163
rect 80 -164 81 -163
rect 81 -164 82 -163
rect 82 -164 83 -163
rect 83 -164 84 -163
rect 84 -164 85 -163
rect 85 -164 86 -163
rect 86 -164 87 -163
rect 87 -164 88 -163
rect 88 -164 89 -163
rect 89 -164 90 -163
rect 90 -164 91 -163
rect 91 -164 92 -163
rect 92 -164 93 -163
rect 93 -164 94 -163
rect 94 -164 95 -163
rect 95 -164 96 -163
rect 96 -164 97 -163
rect 97 -164 98 -163
rect 98 -164 99 -163
rect 99 -164 100 -163
rect 100 -164 101 -163
rect 101 -164 102 -163
rect 102 -164 103 -163
rect 103 -164 104 -163
rect 104 -164 105 -163
rect 105 -164 106 -163
rect 106 -164 107 -163
rect 107 -164 108 -163
rect 108 -164 109 -163
rect 109 -164 110 -163
rect 110 -164 111 -163
rect 111 -164 112 -163
rect 112 -164 113 -163
rect 113 -164 114 -163
rect 114 -164 115 -163
rect 115 -164 116 -163
rect 116 -164 117 -163
rect 117 -164 118 -163
rect 118 -164 119 -163
rect 119 -164 120 -163
rect 120 -164 121 -163
rect 121 -164 122 -163
rect 122 -164 123 -163
rect 123 -164 124 -163
rect 124 -164 125 -163
rect 125 -164 126 -163
rect 126 -164 127 -163
rect 127 -164 128 -163
rect 128 -164 129 -163
rect 129 -164 130 -163
rect 130 -164 131 -163
rect 131 -164 132 -163
rect 132 -164 133 -163
rect 133 -164 134 -163
rect 134 -164 135 -163
rect 135 -164 136 -163
rect 136 -164 137 -163
rect 137 -164 138 -163
rect 138 -164 139 -163
rect 139 -164 140 -163
rect 140 -164 141 -163
rect 141 -164 142 -163
rect 142 -164 143 -163
rect 143 -164 144 -163
rect 144 -164 145 -163
rect 145 -164 146 -163
rect 146 -164 147 -163
rect 147 -164 148 -163
rect 148 -164 149 -163
rect 149 -164 150 -163
rect 150 -164 151 -163
rect 151 -164 152 -163
rect 152 -164 153 -163
rect 153 -164 154 -163
rect 154 -164 155 -163
rect 155 -164 156 -163
rect 156 -164 157 -163
rect 157 -164 158 -163
rect 158 -164 159 -163
rect 159 -164 160 -163
rect 160 -164 161 -163
rect 161 -164 162 -163
rect 162 -164 163 -163
rect 163 -164 164 -163
rect 164 -164 165 -163
rect 165 -164 166 -163
rect 166 -164 167 -163
rect 167 -164 168 -163
rect 168 -164 169 -163
rect 169 -164 170 -163
rect 170 -164 171 -163
rect 171 -164 172 -163
rect 172 -164 173 -163
rect 173 -164 174 -163
rect 174 -164 175 -163
rect 175 -164 176 -163
rect 176 -164 177 -163
rect 177 -164 178 -163
rect 178 -164 179 -163
rect 179 -164 180 -163
rect 180 -164 181 -163
rect 181 -164 182 -163
rect 182 -164 183 -163
rect 183 -164 184 -163
rect 184 -164 185 -163
rect 185 -164 186 -163
rect 186 -164 187 -163
rect 187 -164 188 -163
rect 188 -164 189 -163
rect 189 -164 190 -163
rect 190 -164 191 -163
rect 191 -164 192 -163
rect 192 -164 193 -163
rect 193 -164 194 -163
rect 194 -164 195 -163
rect 195 -164 196 -163
rect 196 -164 197 -163
rect 197 -164 198 -163
rect 198 -164 199 -163
rect 199 -164 200 -163
rect 200 -164 201 -163
rect 201 -164 202 -163
rect 202 -164 203 -163
rect 203 -164 204 -163
rect 204 -164 205 -163
rect 205 -164 206 -163
rect 206 -164 207 -163
rect 207 -164 208 -163
rect 208 -164 209 -163
rect 209 -164 210 -163
rect 210 -164 211 -163
rect 211 -164 212 -163
rect 212 -164 213 -163
rect 213 -164 214 -163
rect 214 -164 215 -163
rect 215 -164 216 -163
rect 216 -164 217 -163
rect 217 -164 218 -163
rect 218 -164 219 -163
rect 219 -164 220 -163
rect 220 -164 221 -163
rect 221 -164 222 -163
rect 222 -164 223 -163
rect 223 -164 224 -163
rect 224 -164 225 -163
rect 225 -164 226 -163
rect 226 -164 227 -163
rect 227 -164 228 -163
rect 228 -164 229 -163
rect 229 -164 230 -163
rect 230 -164 231 -163
rect 231 -164 232 -163
rect 232 -164 233 -163
rect 233 -164 234 -163
rect 234 -164 235 -163
rect 235 -164 236 -163
rect 236 -164 237 -163
rect 237 -164 238 -163
rect 238 -164 239 -163
rect 239 -164 240 -163
rect 240 -164 241 -163
rect 241 -164 242 -163
rect 242 -164 243 -163
rect 243 -164 244 -163
rect 244 -164 245 -163
rect 245 -164 246 -163
rect 246 -164 247 -163
rect 247 -164 248 -163
rect 248 -164 249 -163
rect 249 -164 250 -163
rect 250 -164 251 -163
rect 251 -164 252 -163
rect 252 -164 253 -163
rect 253 -164 254 -163
rect 254 -164 255 -163
rect 255 -164 256 -163
rect 256 -164 257 -163
rect 257 -164 258 -163
rect 258 -164 259 -163
rect 259 -164 260 -163
rect 260 -164 261 -163
rect 261 -164 262 -163
rect 262 -164 263 -163
rect 263 -164 264 -163
rect 264 -164 265 -163
rect 265 -164 266 -163
rect 266 -164 267 -163
rect 267 -164 268 -163
rect 268 -164 269 -163
rect 269 -164 270 -163
rect 270 -164 271 -163
rect 271 -164 272 -163
rect 272 -164 273 -163
rect 273 -164 274 -163
rect 274 -164 275 -163
rect 275 -164 276 -163
rect 276 -164 277 -163
rect 277 -164 278 -163
rect 278 -164 279 -163
rect 279 -164 280 -163
rect 280 -164 281 -163
rect 281 -164 282 -163
rect 282 -164 283 -163
rect 283 -164 284 -163
rect 284 -164 285 -163
rect 285 -164 286 -163
rect 286 -164 287 -163
rect 287 -164 288 -163
rect 288 -164 289 -163
rect 289 -164 290 -163
rect 290 -164 291 -163
rect 291 -164 292 -163
rect 292 -164 293 -163
rect 293 -164 294 -163
rect 294 -164 295 -163
rect 295 -164 296 -163
rect 296 -164 297 -163
rect 297 -164 298 -163
rect 298 -164 299 -163
rect 299 -164 300 -163
rect 300 -164 301 -163
rect 301 -164 302 -163
rect 302 -164 303 -163
rect 303 -164 304 -163
rect 304 -164 305 -163
rect 305 -164 306 -163
rect 306 -164 307 -163
rect 307 -164 308 -163
rect 308 -164 309 -163
rect 309 -164 310 -163
rect 310 -164 311 -163
rect 311 -164 312 -163
rect 312 -164 313 -163
rect 313 -164 314 -163
rect 314 -164 315 -163
rect 315 -164 316 -163
rect 316 -164 317 -163
rect 317 -164 318 -163
rect 318 -164 319 -163
rect 319 -164 320 -163
rect 320 -164 321 -163
rect 321 -164 322 -163
rect 322 -164 323 -163
rect 323 -164 324 -163
rect 324 -164 325 -163
rect 325 -164 326 -163
rect 326 -164 327 -163
rect 327 -164 328 -163
rect 328 -164 329 -163
rect 329 -164 330 -163
rect 330 -164 331 -163
rect 331 -164 332 -163
rect 332 -164 333 -163
rect 333 -164 334 -163
rect 334 -164 335 -163
rect 335 -164 336 -163
rect 336 -164 337 -163
rect 337 -164 338 -163
rect 338 -164 339 -163
rect 339 -164 340 -163
rect 340 -164 341 -163
rect 341 -164 342 -163
rect 342 -164 343 -163
rect 343 -164 344 -163
rect 344 -164 345 -163
rect 345 -164 346 -163
rect 346 -164 347 -163
rect 347 -164 348 -163
rect 348 -164 349 -163
rect 349 -164 350 -163
rect 350 -164 351 -163
rect 351 -164 352 -163
rect 352 -164 353 -163
rect 353 -164 354 -163
rect 354 -164 355 -163
rect 355 -164 356 -163
rect 356 -164 357 -163
rect 357 -164 358 -163
rect 358 -164 359 -163
rect 359 -164 360 -163
rect 360 -164 361 -163
rect 361 -164 362 -163
rect 362 -164 363 -163
rect 363 -164 364 -163
rect 364 -164 365 -163
rect 365 -164 366 -163
rect 366 -164 367 -163
rect 367 -164 368 -163
rect 368 -164 369 -163
rect 369 -164 370 -163
rect 370 -164 371 -163
rect 371 -164 372 -163
rect 372 -164 373 -163
rect 373 -164 374 -163
rect 374 -164 375 -163
rect 375 -164 376 -163
rect 376 -164 377 -163
rect 377 -164 378 -163
rect 378 -164 379 -163
rect 379 -164 380 -163
rect 380 -164 381 -163
rect 381 -164 382 -163
rect 382 -164 383 -163
rect 383 -164 384 -163
rect 384 -164 385 -163
rect 385 -164 386 -163
rect 386 -164 387 -163
rect 387 -164 388 -163
rect 388 -164 389 -163
rect 389 -164 390 -163
rect 390 -164 391 -163
rect 391 -164 392 -163
rect 392 -164 393 -163
rect 393 -164 394 -163
rect 394 -164 395 -163
rect 395 -164 396 -163
rect 396 -164 397 -163
rect 397 -164 398 -163
rect 398 -164 399 -163
rect 399 -164 400 -163
rect 400 -164 401 -163
rect 401 -164 402 -163
rect 402 -164 403 -163
rect 403 -164 404 -163
rect 404 -164 405 -163
rect 405 -164 406 -163
rect 406 -164 407 -163
rect 407 -164 408 -163
rect 408 -164 409 -163
rect 409 -164 410 -163
rect 410 -164 411 -163
rect 411 -164 412 -163
rect 412 -164 413 -163
rect 413 -164 414 -163
rect 414 -164 415 -163
rect 415 -164 416 -163
rect 416 -164 417 -163
rect 417 -164 418 -163
rect 418 -164 419 -163
rect 419 -164 420 -163
rect 420 -164 421 -163
rect 421 -164 422 -163
rect 422 -164 423 -163
rect 423 -164 424 -163
rect 424 -164 425 -163
rect 425 -164 426 -163
rect 426 -164 427 -163
rect 427 -164 428 -163
rect 428 -164 429 -163
rect 429 -164 430 -163
rect 430 -164 431 -163
rect 431 -164 432 -163
rect 432 -164 433 -163
rect 433 -164 434 -163
rect 434 -164 435 -163
rect 435 -164 436 -163
rect 436 -164 437 -163
rect 437 -164 438 -163
rect 438 -164 439 -163
rect 439 -164 440 -163
rect 440 -164 441 -163
rect 441 -164 442 -163
rect 442 -164 443 -163
rect 443 -164 444 -163
rect 444 -164 445 -163
rect 445 -164 446 -163
rect 446 -164 447 -163
rect 447 -164 448 -163
rect 448 -164 449 -163
rect 449 -164 450 -163
rect 450 -164 451 -163
rect 451 -164 452 -163
rect 452 -164 453 -163
rect 453 -164 454 -163
rect 454 -164 455 -163
rect 455 -164 456 -163
rect 456 -164 457 -163
rect 457 -164 458 -163
rect 458 -164 459 -163
rect 459 -164 460 -163
rect 460 -164 461 -163
rect 461 -164 462 -163
rect 462 -164 463 -163
rect 463 -164 464 -163
rect 464 -164 465 -163
rect 465 -164 466 -163
rect 466 -164 467 -163
rect 467 -164 468 -163
rect 468 -164 469 -163
rect 469 -164 470 -163
rect 470 -164 471 -163
rect 471 -164 472 -163
rect 472 -164 473 -163
rect 473 -164 474 -163
rect 474 -164 475 -163
rect 475 -164 476 -163
rect 476 -164 477 -163
rect 477 -164 478 -163
rect 478 -164 479 -163
rect 479 -164 480 -163
rect 2 -165 3 -164
rect 3 -165 4 -164
rect 4 -165 5 -164
rect 5 -165 6 -164
rect 6 -165 7 -164
rect 7 -165 8 -164
rect 8 -165 9 -164
rect 9 -165 10 -164
rect 10 -165 11 -164
rect 11 -165 12 -164
rect 12 -165 13 -164
rect 13 -165 14 -164
rect 14 -165 15 -164
rect 15 -165 16 -164
rect 16 -165 17 -164
rect 17 -165 18 -164
rect 18 -165 19 -164
rect 19 -165 20 -164
rect 20 -165 21 -164
rect 21 -165 22 -164
rect 22 -165 23 -164
rect 23 -165 24 -164
rect 24 -165 25 -164
rect 25 -165 26 -164
rect 26 -165 27 -164
rect 27 -165 28 -164
rect 28 -165 29 -164
rect 29 -165 30 -164
rect 30 -165 31 -164
rect 31 -165 32 -164
rect 32 -165 33 -164
rect 33 -165 34 -164
rect 34 -165 35 -164
rect 35 -165 36 -164
rect 36 -165 37 -164
rect 37 -165 38 -164
rect 38 -165 39 -164
rect 39 -165 40 -164
rect 40 -165 41 -164
rect 41 -165 42 -164
rect 42 -165 43 -164
rect 43 -165 44 -164
rect 44 -165 45 -164
rect 45 -165 46 -164
rect 46 -165 47 -164
rect 47 -165 48 -164
rect 48 -165 49 -164
rect 49 -165 50 -164
rect 50 -165 51 -164
rect 51 -165 52 -164
rect 52 -165 53 -164
rect 53 -165 54 -164
rect 54 -165 55 -164
rect 55 -165 56 -164
rect 56 -165 57 -164
rect 57 -165 58 -164
rect 58 -165 59 -164
rect 59 -165 60 -164
rect 60 -165 61 -164
rect 61 -165 62 -164
rect 62 -165 63 -164
rect 63 -165 64 -164
rect 64 -165 65 -164
rect 65 -165 66 -164
rect 66 -165 67 -164
rect 67 -165 68 -164
rect 68 -165 69 -164
rect 69 -165 70 -164
rect 70 -165 71 -164
rect 71 -165 72 -164
rect 72 -165 73 -164
rect 73 -165 74 -164
rect 74 -165 75 -164
rect 75 -165 76 -164
rect 76 -165 77 -164
rect 77 -165 78 -164
rect 78 -165 79 -164
rect 79 -165 80 -164
rect 80 -165 81 -164
rect 81 -165 82 -164
rect 82 -165 83 -164
rect 83 -165 84 -164
rect 84 -165 85 -164
rect 85 -165 86 -164
rect 86 -165 87 -164
rect 87 -165 88 -164
rect 88 -165 89 -164
rect 89 -165 90 -164
rect 90 -165 91 -164
rect 91 -165 92 -164
rect 92 -165 93 -164
rect 93 -165 94 -164
rect 94 -165 95 -164
rect 95 -165 96 -164
rect 96 -165 97 -164
rect 97 -165 98 -164
rect 98 -165 99 -164
rect 99 -165 100 -164
rect 100 -165 101 -164
rect 101 -165 102 -164
rect 102 -165 103 -164
rect 103 -165 104 -164
rect 104 -165 105 -164
rect 105 -165 106 -164
rect 106 -165 107 -164
rect 107 -165 108 -164
rect 108 -165 109 -164
rect 109 -165 110 -164
rect 110 -165 111 -164
rect 111 -165 112 -164
rect 112 -165 113 -164
rect 113 -165 114 -164
rect 114 -165 115 -164
rect 115 -165 116 -164
rect 116 -165 117 -164
rect 117 -165 118 -164
rect 118 -165 119 -164
rect 119 -165 120 -164
rect 120 -165 121 -164
rect 121 -165 122 -164
rect 122 -165 123 -164
rect 123 -165 124 -164
rect 124 -165 125 -164
rect 125 -165 126 -164
rect 126 -165 127 -164
rect 127 -165 128 -164
rect 128 -165 129 -164
rect 129 -165 130 -164
rect 130 -165 131 -164
rect 131 -165 132 -164
rect 132 -165 133 -164
rect 133 -165 134 -164
rect 134 -165 135 -164
rect 135 -165 136 -164
rect 136 -165 137 -164
rect 137 -165 138 -164
rect 138 -165 139 -164
rect 139 -165 140 -164
rect 140 -165 141 -164
rect 141 -165 142 -164
rect 142 -165 143 -164
rect 143 -165 144 -164
rect 144 -165 145 -164
rect 145 -165 146 -164
rect 146 -165 147 -164
rect 147 -165 148 -164
rect 148 -165 149 -164
rect 149 -165 150 -164
rect 150 -165 151 -164
rect 151 -165 152 -164
rect 152 -165 153 -164
rect 153 -165 154 -164
rect 154 -165 155 -164
rect 155 -165 156 -164
rect 156 -165 157 -164
rect 157 -165 158 -164
rect 158 -165 159 -164
rect 159 -165 160 -164
rect 160 -165 161 -164
rect 161 -165 162 -164
rect 162 -165 163 -164
rect 163 -165 164 -164
rect 164 -165 165 -164
rect 165 -165 166 -164
rect 166 -165 167 -164
rect 167 -165 168 -164
rect 168 -165 169 -164
rect 169 -165 170 -164
rect 170 -165 171 -164
rect 171 -165 172 -164
rect 172 -165 173 -164
rect 173 -165 174 -164
rect 174 -165 175 -164
rect 175 -165 176 -164
rect 176 -165 177 -164
rect 177 -165 178 -164
rect 178 -165 179 -164
rect 179 -165 180 -164
rect 180 -165 181 -164
rect 181 -165 182 -164
rect 182 -165 183 -164
rect 183 -165 184 -164
rect 184 -165 185 -164
rect 185 -165 186 -164
rect 186 -165 187 -164
rect 187 -165 188 -164
rect 188 -165 189 -164
rect 189 -165 190 -164
rect 190 -165 191 -164
rect 191 -165 192 -164
rect 192 -165 193 -164
rect 193 -165 194 -164
rect 194 -165 195 -164
rect 195 -165 196 -164
rect 196 -165 197 -164
rect 197 -165 198 -164
rect 198 -165 199 -164
rect 199 -165 200 -164
rect 200 -165 201 -164
rect 201 -165 202 -164
rect 202 -165 203 -164
rect 203 -165 204 -164
rect 204 -165 205 -164
rect 205 -165 206 -164
rect 206 -165 207 -164
rect 207 -165 208 -164
rect 208 -165 209 -164
rect 209 -165 210 -164
rect 210 -165 211 -164
rect 211 -165 212 -164
rect 212 -165 213 -164
rect 213 -165 214 -164
rect 214 -165 215 -164
rect 215 -165 216 -164
rect 216 -165 217 -164
rect 217 -165 218 -164
rect 218 -165 219 -164
rect 219 -165 220 -164
rect 220 -165 221 -164
rect 221 -165 222 -164
rect 222 -165 223 -164
rect 223 -165 224 -164
rect 224 -165 225 -164
rect 225 -165 226 -164
rect 226 -165 227 -164
rect 227 -165 228 -164
rect 228 -165 229 -164
rect 229 -165 230 -164
rect 230 -165 231 -164
rect 231 -165 232 -164
rect 232 -165 233 -164
rect 233 -165 234 -164
rect 234 -165 235 -164
rect 235 -165 236 -164
rect 236 -165 237 -164
rect 237 -165 238 -164
rect 238 -165 239 -164
rect 239 -165 240 -164
rect 240 -165 241 -164
rect 241 -165 242 -164
rect 242 -165 243 -164
rect 243 -165 244 -164
rect 244 -165 245 -164
rect 245 -165 246 -164
rect 246 -165 247 -164
rect 247 -165 248 -164
rect 248 -165 249 -164
rect 249 -165 250 -164
rect 250 -165 251 -164
rect 251 -165 252 -164
rect 252 -165 253 -164
rect 253 -165 254 -164
rect 254 -165 255 -164
rect 255 -165 256 -164
rect 256 -165 257 -164
rect 257 -165 258 -164
rect 258 -165 259 -164
rect 259 -165 260 -164
rect 260 -165 261 -164
rect 261 -165 262 -164
rect 262 -165 263 -164
rect 263 -165 264 -164
rect 264 -165 265 -164
rect 265 -165 266 -164
rect 266 -165 267 -164
rect 267 -165 268 -164
rect 268 -165 269 -164
rect 269 -165 270 -164
rect 270 -165 271 -164
rect 271 -165 272 -164
rect 272 -165 273 -164
rect 273 -165 274 -164
rect 274 -165 275 -164
rect 275 -165 276 -164
rect 276 -165 277 -164
rect 277 -165 278 -164
rect 278 -165 279 -164
rect 279 -165 280 -164
rect 280 -165 281 -164
rect 281 -165 282 -164
rect 282 -165 283 -164
rect 283 -165 284 -164
rect 284 -165 285 -164
rect 285 -165 286 -164
rect 286 -165 287 -164
rect 287 -165 288 -164
rect 288 -165 289 -164
rect 289 -165 290 -164
rect 290 -165 291 -164
rect 291 -165 292 -164
rect 292 -165 293 -164
rect 293 -165 294 -164
rect 294 -165 295 -164
rect 295 -165 296 -164
rect 296 -165 297 -164
rect 297 -165 298 -164
rect 298 -165 299 -164
rect 299 -165 300 -164
rect 300 -165 301 -164
rect 301 -165 302 -164
rect 302 -165 303 -164
rect 303 -165 304 -164
rect 304 -165 305 -164
rect 305 -165 306 -164
rect 306 -165 307 -164
rect 307 -165 308 -164
rect 308 -165 309 -164
rect 309 -165 310 -164
rect 310 -165 311 -164
rect 311 -165 312 -164
rect 312 -165 313 -164
rect 313 -165 314 -164
rect 314 -165 315 -164
rect 315 -165 316 -164
rect 316 -165 317 -164
rect 317 -165 318 -164
rect 318 -165 319 -164
rect 319 -165 320 -164
rect 320 -165 321 -164
rect 321 -165 322 -164
rect 322 -165 323 -164
rect 323 -165 324 -164
rect 324 -165 325 -164
rect 325 -165 326 -164
rect 326 -165 327 -164
rect 327 -165 328 -164
rect 328 -165 329 -164
rect 329 -165 330 -164
rect 330 -165 331 -164
rect 331 -165 332 -164
rect 332 -165 333 -164
rect 333 -165 334 -164
rect 334 -165 335 -164
rect 335 -165 336 -164
rect 336 -165 337 -164
rect 337 -165 338 -164
rect 338 -165 339 -164
rect 339 -165 340 -164
rect 340 -165 341 -164
rect 341 -165 342 -164
rect 342 -165 343 -164
rect 343 -165 344 -164
rect 344 -165 345 -164
rect 345 -165 346 -164
rect 346 -165 347 -164
rect 347 -165 348 -164
rect 348 -165 349 -164
rect 349 -165 350 -164
rect 350 -165 351 -164
rect 351 -165 352 -164
rect 352 -165 353 -164
rect 353 -165 354 -164
rect 354 -165 355 -164
rect 355 -165 356 -164
rect 356 -165 357 -164
rect 357 -165 358 -164
rect 358 -165 359 -164
rect 359 -165 360 -164
rect 360 -165 361 -164
rect 361 -165 362 -164
rect 362 -165 363 -164
rect 363 -165 364 -164
rect 364 -165 365 -164
rect 365 -165 366 -164
rect 366 -165 367 -164
rect 367 -165 368 -164
rect 368 -165 369 -164
rect 369 -165 370 -164
rect 370 -165 371 -164
rect 371 -165 372 -164
rect 372 -165 373 -164
rect 373 -165 374 -164
rect 374 -165 375 -164
rect 375 -165 376 -164
rect 376 -165 377 -164
rect 377 -165 378 -164
rect 378 -165 379 -164
rect 379 -165 380 -164
rect 380 -165 381 -164
rect 381 -165 382 -164
rect 382 -165 383 -164
rect 383 -165 384 -164
rect 384 -165 385 -164
rect 385 -165 386 -164
rect 386 -165 387 -164
rect 387 -165 388 -164
rect 388 -165 389 -164
rect 389 -165 390 -164
rect 390 -165 391 -164
rect 391 -165 392 -164
rect 392 -165 393 -164
rect 393 -165 394 -164
rect 394 -165 395 -164
rect 395 -165 396 -164
rect 396 -165 397 -164
rect 397 -165 398 -164
rect 398 -165 399 -164
rect 399 -165 400 -164
rect 400 -165 401 -164
rect 401 -165 402 -164
rect 402 -165 403 -164
rect 403 -165 404 -164
rect 404 -165 405 -164
rect 405 -165 406 -164
rect 406 -165 407 -164
rect 407 -165 408 -164
rect 408 -165 409 -164
rect 409 -165 410 -164
rect 410 -165 411 -164
rect 411 -165 412 -164
rect 412 -165 413 -164
rect 413 -165 414 -164
rect 414 -165 415 -164
rect 415 -165 416 -164
rect 416 -165 417 -164
rect 417 -165 418 -164
rect 418 -165 419 -164
rect 419 -165 420 -164
rect 420 -165 421 -164
rect 421 -165 422 -164
rect 422 -165 423 -164
rect 423 -165 424 -164
rect 424 -165 425 -164
rect 425 -165 426 -164
rect 426 -165 427 -164
rect 427 -165 428 -164
rect 428 -165 429 -164
rect 429 -165 430 -164
rect 430 -165 431 -164
rect 431 -165 432 -164
rect 432 -165 433 -164
rect 433 -165 434 -164
rect 434 -165 435 -164
rect 435 -165 436 -164
rect 436 -165 437 -164
rect 437 -165 438 -164
rect 438 -165 439 -164
rect 439 -165 440 -164
rect 440 -165 441 -164
rect 441 -165 442 -164
rect 442 -165 443 -164
rect 443 -165 444 -164
rect 444 -165 445 -164
rect 445 -165 446 -164
rect 446 -165 447 -164
rect 447 -165 448 -164
rect 448 -165 449 -164
rect 449 -165 450 -164
rect 450 -165 451 -164
rect 451 -165 452 -164
rect 452 -165 453 -164
rect 453 -165 454 -164
rect 454 -165 455 -164
rect 455 -165 456 -164
rect 456 -165 457 -164
rect 457 -165 458 -164
rect 458 -165 459 -164
rect 459 -165 460 -164
rect 460 -165 461 -164
rect 461 -165 462 -164
rect 462 -165 463 -164
rect 463 -165 464 -164
rect 464 -165 465 -164
rect 465 -165 466 -164
rect 466 -165 467 -164
rect 467 -165 468 -164
rect 468 -165 469 -164
rect 469 -165 470 -164
rect 470 -165 471 -164
rect 471 -165 472 -164
rect 472 -165 473 -164
rect 473 -165 474 -164
rect 474 -165 475 -164
rect 475 -165 476 -164
rect 476 -165 477 -164
rect 477 -165 478 -164
rect 478 -165 479 -164
rect 479 -165 480 -164
rect 2 -166 3 -165
rect 3 -166 4 -165
rect 4 -166 5 -165
rect 5 -166 6 -165
rect 6 -166 7 -165
rect 7 -166 8 -165
rect 8 -166 9 -165
rect 9 -166 10 -165
rect 10 -166 11 -165
rect 11 -166 12 -165
rect 12 -166 13 -165
rect 13 -166 14 -165
rect 14 -166 15 -165
rect 15 -166 16 -165
rect 16 -166 17 -165
rect 17 -166 18 -165
rect 18 -166 19 -165
rect 19 -166 20 -165
rect 20 -166 21 -165
rect 21 -166 22 -165
rect 22 -166 23 -165
rect 23 -166 24 -165
rect 24 -166 25 -165
rect 25 -166 26 -165
rect 26 -166 27 -165
rect 27 -166 28 -165
rect 28 -166 29 -165
rect 29 -166 30 -165
rect 30 -166 31 -165
rect 31 -166 32 -165
rect 32 -166 33 -165
rect 33 -166 34 -165
rect 34 -166 35 -165
rect 35 -166 36 -165
rect 36 -166 37 -165
rect 37 -166 38 -165
rect 38 -166 39 -165
rect 39 -166 40 -165
rect 40 -166 41 -165
rect 41 -166 42 -165
rect 42 -166 43 -165
rect 43 -166 44 -165
rect 44 -166 45 -165
rect 45 -166 46 -165
rect 46 -166 47 -165
rect 47 -166 48 -165
rect 48 -166 49 -165
rect 49 -166 50 -165
rect 50 -166 51 -165
rect 51 -166 52 -165
rect 52 -166 53 -165
rect 53 -166 54 -165
rect 54 -166 55 -165
rect 55 -166 56 -165
rect 56 -166 57 -165
rect 57 -166 58 -165
rect 58 -166 59 -165
rect 59 -166 60 -165
rect 60 -166 61 -165
rect 61 -166 62 -165
rect 62 -166 63 -165
rect 63 -166 64 -165
rect 64 -166 65 -165
rect 65 -166 66 -165
rect 66 -166 67 -165
rect 67 -166 68 -165
rect 68 -166 69 -165
rect 69 -166 70 -165
rect 70 -166 71 -165
rect 71 -166 72 -165
rect 72 -166 73 -165
rect 73 -166 74 -165
rect 74 -166 75 -165
rect 75 -166 76 -165
rect 76 -166 77 -165
rect 77 -166 78 -165
rect 78 -166 79 -165
rect 79 -166 80 -165
rect 80 -166 81 -165
rect 81 -166 82 -165
rect 82 -166 83 -165
rect 83 -166 84 -165
rect 84 -166 85 -165
rect 85 -166 86 -165
rect 86 -166 87 -165
rect 87 -166 88 -165
rect 88 -166 89 -165
rect 89 -166 90 -165
rect 90 -166 91 -165
rect 91 -166 92 -165
rect 92 -166 93 -165
rect 93 -166 94 -165
rect 94 -166 95 -165
rect 95 -166 96 -165
rect 96 -166 97 -165
rect 97 -166 98 -165
rect 98 -166 99 -165
rect 99 -166 100 -165
rect 100 -166 101 -165
rect 101 -166 102 -165
rect 102 -166 103 -165
rect 103 -166 104 -165
rect 104 -166 105 -165
rect 105 -166 106 -165
rect 106 -166 107 -165
rect 107 -166 108 -165
rect 108 -166 109 -165
rect 109 -166 110 -165
rect 110 -166 111 -165
rect 111 -166 112 -165
rect 112 -166 113 -165
rect 113 -166 114 -165
rect 114 -166 115 -165
rect 115 -166 116 -165
rect 116 -166 117 -165
rect 117 -166 118 -165
rect 118 -166 119 -165
rect 119 -166 120 -165
rect 120 -166 121 -165
rect 121 -166 122 -165
rect 122 -166 123 -165
rect 123 -166 124 -165
rect 124 -166 125 -165
rect 125 -166 126 -165
rect 126 -166 127 -165
rect 127 -166 128 -165
rect 128 -166 129 -165
rect 129 -166 130 -165
rect 130 -166 131 -165
rect 131 -166 132 -165
rect 132 -166 133 -165
rect 133 -166 134 -165
rect 134 -166 135 -165
rect 135 -166 136 -165
rect 136 -166 137 -165
rect 137 -166 138 -165
rect 138 -166 139 -165
rect 139 -166 140 -165
rect 140 -166 141 -165
rect 141 -166 142 -165
rect 142 -166 143 -165
rect 143 -166 144 -165
rect 144 -166 145 -165
rect 145 -166 146 -165
rect 146 -166 147 -165
rect 147 -166 148 -165
rect 148 -166 149 -165
rect 149 -166 150 -165
rect 150 -166 151 -165
rect 151 -166 152 -165
rect 152 -166 153 -165
rect 153 -166 154 -165
rect 154 -166 155 -165
rect 155 -166 156 -165
rect 156 -166 157 -165
rect 157 -166 158 -165
rect 158 -166 159 -165
rect 159 -166 160 -165
rect 160 -166 161 -165
rect 161 -166 162 -165
rect 162 -166 163 -165
rect 163 -166 164 -165
rect 164 -166 165 -165
rect 165 -166 166 -165
rect 166 -166 167 -165
rect 167 -166 168 -165
rect 168 -166 169 -165
rect 169 -166 170 -165
rect 170 -166 171 -165
rect 171 -166 172 -165
rect 172 -166 173 -165
rect 173 -166 174 -165
rect 174 -166 175 -165
rect 175 -166 176 -165
rect 176 -166 177 -165
rect 177 -166 178 -165
rect 178 -166 179 -165
rect 179 -166 180 -165
rect 180 -166 181 -165
rect 181 -166 182 -165
rect 182 -166 183 -165
rect 183 -166 184 -165
rect 184 -166 185 -165
rect 185 -166 186 -165
rect 186 -166 187 -165
rect 187 -166 188 -165
rect 188 -166 189 -165
rect 189 -166 190 -165
rect 190 -166 191 -165
rect 191 -166 192 -165
rect 192 -166 193 -165
rect 193 -166 194 -165
rect 194 -166 195 -165
rect 195 -166 196 -165
rect 196 -166 197 -165
rect 197 -166 198 -165
rect 198 -166 199 -165
rect 199 -166 200 -165
rect 200 -166 201 -165
rect 201 -166 202 -165
rect 202 -166 203 -165
rect 203 -166 204 -165
rect 204 -166 205 -165
rect 205 -166 206 -165
rect 206 -166 207 -165
rect 207 -166 208 -165
rect 208 -166 209 -165
rect 209 -166 210 -165
rect 210 -166 211 -165
rect 211 -166 212 -165
rect 212 -166 213 -165
rect 213 -166 214 -165
rect 214 -166 215 -165
rect 215 -166 216 -165
rect 216 -166 217 -165
rect 217 -166 218 -165
rect 218 -166 219 -165
rect 219 -166 220 -165
rect 220 -166 221 -165
rect 221 -166 222 -165
rect 222 -166 223 -165
rect 223 -166 224 -165
rect 224 -166 225 -165
rect 225 -166 226 -165
rect 226 -166 227 -165
rect 227 -166 228 -165
rect 228 -166 229 -165
rect 229 -166 230 -165
rect 230 -166 231 -165
rect 231 -166 232 -165
rect 232 -166 233 -165
rect 233 -166 234 -165
rect 234 -166 235 -165
rect 235 -166 236 -165
rect 236 -166 237 -165
rect 237 -166 238 -165
rect 238 -166 239 -165
rect 239 -166 240 -165
rect 240 -166 241 -165
rect 241 -166 242 -165
rect 242 -166 243 -165
rect 243 -166 244 -165
rect 244 -166 245 -165
rect 245 -166 246 -165
rect 246 -166 247 -165
rect 247 -166 248 -165
rect 248 -166 249 -165
rect 249 -166 250 -165
rect 250 -166 251 -165
rect 251 -166 252 -165
rect 252 -166 253 -165
rect 253 -166 254 -165
rect 254 -166 255 -165
rect 255 -166 256 -165
rect 256 -166 257 -165
rect 257 -166 258 -165
rect 258 -166 259 -165
rect 259 -166 260 -165
rect 260 -166 261 -165
rect 261 -166 262 -165
rect 262 -166 263 -165
rect 263 -166 264 -165
rect 264 -166 265 -165
rect 265 -166 266 -165
rect 266 -166 267 -165
rect 267 -166 268 -165
rect 268 -166 269 -165
rect 269 -166 270 -165
rect 270 -166 271 -165
rect 271 -166 272 -165
rect 272 -166 273 -165
rect 273 -166 274 -165
rect 274 -166 275 -165
rect 275 -166 276 -165
rect 276 -166 277 -165
rect 277 -166 278 -165
rect 278 -166 279 -165
rect 279 -166 280 -165
rect 280 -166 281 -165
rect 281 -166 282 -165
rect 282 -166 283 -165
rect 283 -166 284 -165
rect 284 -166 285 -165
rect 285 -166 286 -165
rect 286 -166 287 -165
rect 287 -166 288 -165
rect 288 -166 289 -165
rect 289 -166 290 -165
rect 290 -166 291 -165
rect 291 -166 292 -165
rect 292 -166 293 -165
rect 293 -166 294 -165
rect 294 -166 295 -165
rect 295 -166 296 -165
rect 296 -166 297 -165
rect 297 -166 298 -165
rect 298 -166 299 -165
rect 299 -166 300 -165
rect 300 -166 301 -165
rect 301 -166 302 -165
rect 302 -166 303 -165
rect 303 -166 304 -165
rect 304 -166 305 -165
rect 305 -166 306 -165
rect 306 -166 307 -165
rect 307 -166 308 -165
rect 308 -166 309 -165
rect 309 -166 310 -165
rect 310 -166 311 -165
rect 311 -166 312 -165
rect 312 -166 313 -165
rect 313 -166 314 -165
rect 314 -166 315 -165
rect 315 -166 316 -165
rect 316 -166 317 -165
rect 317 -166 318 -165
rect 318 -166 319 -165
rect 319 -166 320 -165
rect 320 -166 321 -165
rect 321 -166 322 -165
rect 322 -166 323 -165
rect 323 -166 324 -165
rect 324 -166 325 -165
rect 325 -166 326 -165
rect 326 -166 327 -165
rect 327 -166 328 -165
rect 328 -166 329 -165
rect 329 -166 330 -165
rect 330 -166 331 -165
rect 331 -166 332 -165
rect 332 -166 333 -165
rect 333 -166 334 -165
rect 334 -166 335 -165
rect 335 -166 336 -165
rect 336 -166 337 -165
rect 337 -166 338 -165
rect 338 -166 339 -165
rect 339 -166 340 -165
rect 340 -166 341 -165
rect 341 -166 342 -165
rect 342 -166 343 -165
rect 343 -166 344 -165
rect 344 -166 345 -165
rect 345 -166 346 -165
rect 346 -166 347 -165
rect 347 -166 348 -165
rect 348 -166 349 -165
rect 349 -166 350 -165
rect 350 -166 351 -165
rect 351 -166 352 -165
rect 352 -166 353 -165
rect 353 -166 354 -165
rect 354 -166 355 -165
rect 355 -166 356 -165
rect 356 -166 357 -165
rect 357 -166 358 -165
rect 358 -166 359 -165
rect 359 -166 360 -165
rect 360 -166 361 -165
rect 361 -166 362 -165
rect 362 -166 363 -165
rect 363 -166 364 -165
rect 364 -166 365 -165
rect 365 -166 366 -165
rect 366 -166 367 -165
rect 367 -166 368 -165
rect 368 -166 369 -165
rect 369 -166 370 -165
rect 370 -166 371 -165
rect 371 -166 372 -165
rect 372 -166 373 -165
rect 373 -166 374 -165
rect 374 -166 375 -165
rect 375 -166 376 -165
rect 376 -166 377 -165
rect 377 -166 378 -165
rect 378 -166 379 -165
rect 379 -166 380 -165
rect 380 -166 381 -165
rect 381 -166 382 -165
rect 382 -166 383 -165
rect 383 -166 384 -165
rect 384 -166 385 -165
rect 385 -166 386 -165
rect 386 -166 387 -165
rect 387 -166 388 -165
rect 388 -166 389 -165
rect 389 -166 390 -165
rect 390 -166 391 -165
rect 391 -166 392 -165
rect 392 -166 393 -165
rect 393 -166 394 -165
rect 394 -166 395 -165
rect 395 -166 396 -165
rect 396 -166 397 -165
rect 397 -166 398 -165
rect 398 -166 399 -165
rect 399 -166 400 -165
rect 400 -166 401 -165
rect 401 -166 402 -165
rect 402 -166 403 -165
rect 403 -166 404 -165
rect 404 -166 405 -165
rect 405 -166 406 -165
rect 406 -166 407 -165
rect 407 -166 408 -165
rect 408 -166 409 -165
rect 409 -166 410 -165
rect 410 -166 411 -165
rect 411 -166 412 -165
rect 412 -166 413 -165
rect 413 -166 414 -165
rect 414 -166 415 -165
rect 415 -166 416 -165
rect 416 -166 417 -165
rect 417 -166 418 -165
rect 418 -166 419 -165
rect 419 -166 420 -165
rect 420 -166 421 -165
rect 421 -166 422 -165
rect 422 -166 423 -165
rect 423 -166 424 -165
rect 424 -166 425 -165
rect 425 -166 426 -165
rect 426 -166 427 -165
rect 427 -166 428 -165
rect 428 -166 429 -165
rect 429 -166 430 -165
rect 430 -166 431 -165
rect 431 -166 432 -165
rect 432 -166 433 -165
rect 433 -166 434 -165
rect 434 -166 435 -165
rect 435 -166 436 -165
rect 436 -166 437 -165
rect 437 -166 438 -165
rect 438 -166 439 -165
rect 439 -166 440 -165
rect 440 -166 441 -165
rect 441 -166 442 -165
rect 442 -166 443 -165
rect 443 -166 444 -165
rect 444 -166 445 -165
rect 445 -166 446 -165
rect 446 -166 447 -165
rect 447 -166 448 -165
rect 448 -166 449 -165
rect 449 -166 450 -165
rect 450 -166 451 -165
rect 451 -166 452 -165
rect 452 -166 453 -165
rect 453 -166 454 -165
rect 454 -166 455 -165
rect 455 -166 456 -165
rect 456 -166 457 -165
rect 457 -166 458 -165
rect 458 -166 459 -165
rect 459 -166 460 -165
rect 460 -166 461 -165
rect 461 -166 462 -165
rect 462 -166 463 -165
rect 463 -166 464 -165
rect 464 -166 465 -165
rect 465 -166 466 -165
rect 466 -166 467 -165
rect 467 -166 468 -165
rect 468 -166 469 -165
rect 469 -166 470 -165
rect 470 -166 471 -165
rect 471 -166 472 -165
rect 472 -166 473 -165
rect 473 -166 474 -165
rect 474 -166 475 -165
rect 475 -166 476 -165
rect 476 -166 477 -165
rect 477 -166 478 -165
rect 478 -166 479 -165
rect 479 -166 480 -165
rect 2 -167 3 -166
rect 3 -167 4 -166
rect 4 -167 5 -166
rect 5 -167 6 -166
rect 6 -167 7 -166
rect 7 -167 8 -166
rect 8 -167 9 -166
rect 9 -167 10 -166
rect 10 -167 11 -166
rect 11 -167 12 -166
rect 12 -167 13 -166
rect 13 -167 14 -166
rect 14 -167 15 -166
rect 15 -167 16 -166
rect 16 -167 17 -166
rect 17 -167 18 -166
rect 18 -167 19 -166
rect 19 -167 20 -166
rect 20 -167 21 -166
rect 21 -167 22 -166
rect 22 -167 23 -166
rect 23 -167 24 -166
rect 24 -167 25 -166
rect 25 -167 26 -166
rect 26 -167 27 -166
rect 27 -167 28 -166
rect 28 -167 29 -166
rect 29 -167 30 -166
rect 30 -167 31 -166
rect 31 -167 32 -166
rect 32 -167 33 -166
rect 33 -167 34 -166
rect 34 -167 35 -166
rect 35 -167 36 -166
rect 36 -167 37 -166
rect 37 -167 38 -166
rect 38 -167 39 -166
rect 39 -167 40 -166
rect 40 -167 41 -166
rect 41 -167 42 -166
rect 42 -167 43 -166
rect 43 -167 44 -166
rect 44 -167 45 -166
rect 45 -167 46 -166
rect 46 -167 47 -166
rect 47 -167 48 -166
rect 48 -167 49 -166
rect 49 -167 50 -166
rect 50 -167 51 -166
rect 51 -167 52 -166
rect 52 -167 53 -166
rect 53 -167 54 -166
rect 54 -167 55 -166
rect 55 -167 56 -166
rect 56 -167 57 -166
rect 57 -167 58 -166
rect 58 -167 59 -166
rect 59 -167 60 -166
rect 60 -167 61 -166
rect 61 -167 62 -166
rect 62 -167 63 -166
rect 63 -167 64 -166
rect 64 -167 65 -166
rect 65 -167 66 -166
rect 66 -167 67 -166
rect 67 -167 68 -166
rect 68 -167 69 -166
rect 69 -167 70 -166
rect 70 -167 71 -166
rect 71 -167 72 -166
rect 72 -167 73 -166
rect 73 -167 74 -166
rect 74 -167 75 -166
rect 75 -167 76 -166
rect 76 -167 77 -166
rect 77 -167 78 -166
rect 78 -167 79 -166
rect 79 -167 80 -166
rect 80 -167 81 -166
rect 81 -167 82 -166
rect 82 -167 83 -166
rect 83 -167 84 -166
rect 84 -167 85 -166
rect 85 -167 86 -166
rect 86 -167 87 -166
rect 87 -167 88 -166
rect 88 -167 89 -166
rect 89 -167 90 -166
rect 90 -167 91 -166
rect 91 -167 92 -166
rect 92 -167 93 -166
rect 93 -167 94 -166
rect 94 -167 95 -166
rect 95 -167 96 -166
rect 96 -167 97 -166
rect 97 -167 98 -166
rect 98 -167 99 -166
rect 99 -167 100 -166
rect 100 -167 101 -166
rect 101 -167 102 -166
rect 102 -167 103 -166
rect 103 -167 104 -166
rect 104 -167 105 -166
rect 105 -167 106 -166
rect 106 -167 107 -166
rect 107 -167 108 -166
rect 108 -167 109 -166
rect 109 -167 110 -166
rect 110 -167 111 -166
rect 111 -167 112 -166
rect 112 -167 113 -166
rect 113 -167 114 -166
rect 114 -167 115 -166
rect 115 -167 116 -166
rect 116 -167 117 -166
rect 117 -167 118 -166
rect 118 -167 119 -166
rect 119 -167 120 -166
rect 120 -167 121 -166
rect 121 -167 122 -166
rect 122 -167 123 -166
rect 123 -167 124 -166
rect 124 -167 125 -166
rect 125 -167 126 -166
rect 126 -167 127 -166
rect 127 -167 128 -166
rect 128 -167 129 -166
rect 129 -167 130 -166
rect 130 -167 131 -166
rect 131 -167 132 -166
rect 132 -167 133 -166
rect 133 -167 134 -166
rect 134 -167 135 -166
rect 135 -167 136 -166
rect 136 -167 137 -166
rect 137 -167 138 -166
rect 138 -167 139 -166
rect 139 -167 140 -166
rect 140 -167 141 -166
rect 141 -167 142 -166
rect 142 -167 143 -166
rect 143 -167 144 -166
rect 144 -167 145 -166
rect 145 -167 146 -166
rect 146 -167 147 -166
rect 147 -167 148 -166
rect 148 -167 149 -166
rect 149 -167 150 -166
rect 150 -167 151 -166
rect 151 -167 152 -166
rect 152 -167 153 -166
rect 153 -167 154 -166
rect 154 -167 155 -166
rect 155 -167 156 -166
rect 156 -167 157 -166
rect 157 -167 158 -166
rect 158 -167 159 -166
rect 159 -167 160 -166
rect 160 -167 161 -166
rect 161 -167 162 -166
rect 162 -167 163 -166
rect 163 -167 164 -166
rect 164 -167 165 -166
rect 165 -167 166 -166
rect 166 -167 167 -166
rect 167 -167 168 -166
rect 168 -167 169 -166
rect 169 -167 170 -166
rect 170 -167 171 -166
rect 171 -167 172 -166
rect 172 -167 173 -166
rect 173 -167 174 -166
rect 174 -167 175 -166
rect 175 -167 176 -166
rect 176 -167 177 -166
rect 177 -167 178 -166
rect 178 -167 179 -166
rect 179 -167 180 -166
rect 180 -167 181 -166
rect 181 -167 182 -166
rect 182 -167 183 -166
rect 183 -167 184 -166
rect 184 -167 185 -166
rect 185 -167 186 -166
rect 186 -167 187 -166
rect 187 -167 188 -166
rect 188 -167 189 -166
rect 189 -167 190 -166
rect 190 -167 191 -166
rect 191 -167 192 -166
rect 192 -167 193 -166
rect 193 -167 194 -166
rect 194 -167 195 -166
rect 195 -167 196 -166
rect 196 -167 197 -166
rect 197 -167 198 -166
rect 198 -167 199 -166
rect 199 -167 200 -166
rect 200 -167 201 -166
rect 201 -167 202 -166
rect 202 -167 203 -166
rect 203 -167 204 -166
rect 204 -167 205 -166
rect 205 -167 206 -166
rect 206 -167 207 -166
rect 207 -167 208 -166
rect 208 -167 209 -166
rect 209 -167 210 -166
rect 210 -167 211 -166
rect 211 -167 212 -166
rect 212 -167 213 -166
rect 213 -167 214 -166
rect 214 -167 215 -166
rect 215 -167 216 -166
rect 216 -167 217 -166
rect 217 -167 218 -166
rect 218 -167 219 -166
rect 219 -167 220 -166
rect 220 -167 221 -166
rect 221 -167 222 -166
rect 222 -167 223 -166
rect 223 -167 224 -166
rect 224 -167 225 -166
rect 225 -167 226 -166
rect 226 -167 227 -166
rect 227 -167 228 -166
rect 228 -167 229 -166
rect 229 -167 230 -166
rect 230 -167 231 -166
rect 231 -167 232 -166
rect 232 -167 233 -166
rect 233 -167 234 -166
rect 234 -167 235 -166
rect 235 -167 236 -166
rect 236 -167 237 -166
rect 237 -167 238 -166
rect 238 -167 239 -166
rect 239 -167 240 -166
rect 240 -167 241 -166
rect 241 -167 242 -166
rect 242 -167 243 -166
rect 243 -167 244 -166
rect 244 -167 245 -166
rect 245 -167 246 -166
rect 246 -167 247 -166
rect 247 -167 248 -166
rect 248 -167 249 -166
rect 249 -167 250 -166
rect 250 -167 251 -166
rect 251 -167 252 -166
rect 252 -167 253 -166
rect 253 -167 254 -166
rect 254 -167 255 -166
rect 255 -167 256 -166
rect 256 -167 257 -166
rect 257 -167 258 -166
rect 258 -167 259 -166
rect 259 -167 260 -166
rect 260 -167 261 -166
rect 261 -167 262 -166
rect 262 -167 263 -166
rect 263 -167 264 -166
rect 264 -167 265 -166
rect 265 -167 266 -166
rect 266 -167 267 -166
rect 267 -167 268 -166
rect 268 -167 269 -166
rect 269 -167 270 -166
rect 270 -167 271 -166
rect 271 -167 272 -166
rect 272 -167 273 -166
rect 273 -167 274 -166
rect 274 -167 275 -166
rect 275 -167 276 -166
rect 276 -167 277 -166
rect 277 -167 278 -166
rect 278 -167 279 -166
rect 279 -167 280 -166
rect 280 -167 281 -166
rect 281 -167 282 -166
rect 282 -167 283 -166
rect 283 -167 284 -166
rect 284 -167 285 -166
rect 285 -167 286 -166
rect 286 -167 287 -166
rect 287 -167 288 -166
rect 288 -167 289 -166
rect 289 -167 290 -166
rect 290 -167 291 -166
rect 291 -167 292 -166
rect 292 -167 293 -166
rect 293 -167 294 -166
rect 294 -167 295 -166
rect 295 -167 296 -166
rect 296 -167 297 -166
rect 297 -167 298 -166
rect 298 -167 299 -166
rect 299 -167 300 -166
rect 300 -167 301 -166
rect 301 -167 302 -166
rect 302 -167 303 -166
rect 303 -167 304 -166
rect 304 -167 305 -166
rect 305 -167 306 -166
rect 306 -167 307 -166
rect 307 -167 308 -166
rect 308 -167 309 -166
rect 309 -167 310 -166
rect 310 -167 311 -166
rect 311 -167 312 -166
rect 312 -167 313 -166
rect 313 -167 314 -166
rect 314 -167 315 -166
rect 315 -167 316 -166
rect 316 -167 317 -166
rect 317 -167 318 -166
rect 318 -167 319 -166
rect 319 -167 320 -166
rect 320 -167 321 -166
rect 321 -167 322 -166
rect 322 -167 323 -166
rect 323 -167 324 -166
rect 324 -167 325 -166
rect 325 -167 326 -166
rect 326 -167 327 -166
rect 327 -167 328 -166
rect 328 -167 329 -166
rect 329 -167 330 -166
rect 330 -167 331 -166
rect 331 -167 332 -166
rect 332 -167 333 -166
rect 333 -167 334 -166
rect 334 -167 335 -166
rect 335 -167 336 -166
rect 336 -167 337 -166
rect 337 -167 338 -166
rect 338 -167 339 -166
rect 339 -167 340 -166
rect 340 -167 341 -166
rect 341 -167 342 -166
rect 342 -167 343 -166
rect 343 -167 344 -166
rect 344 -167 345 -166
rect 345 -167 346 -166
rect 346 -167 347 -166
rect 347 -167 348 -166
rect 348 -167 349 -166
rect 349 -167 350 -166
rect 350 -167 351 -166
rect 351 -167 352 -166
rect 352 -167 353 -166
rect 353 -167 354 -166
rect 354 -167 355 -166
rect 355 -167 356 -166
rect 356 -167 357 -166
rect 357 -167 358 -166
rect 358 -167 359 -166
rect 359 -167 360 -166
rect 360 -167 361 -166
rect 361 -167 362 -166
rect 362 -167 363 -166
rect 363 -167 364 -166
rect 364 -167 365 -166
rect 365 -167 366 -166
rect 366 -167 367 -166
rect 367 -167 368 -166
rect 368 -167 369 -166
rect 369 -167 370 -166
rect 370 -167 371 -166
rect 371 -167 372 -166
rect 372 -167 373 -166
rect 373 -167 374 -166
rect 374 -167 375 -166
rect 375 -167 376 -166
rect 376 -167 377 -166
rect 377 -167 378 -166
rect 378 -167 379 -166
rect 379 -167 380 -166
rect 380 -167 381 -166
rect 381 -167 382 -166
rect 382 -167 383 -166
rect 383 -167 384 -166
rect 384 -167 385 -166
rect 385 -167 386 -166
rect 386 -167 387 -166
rect 387 -167 388 -166
rect 388 -167 389 -166
rect 389 -167 390 -166
rect 390 -167 391 -166
rect 391 -167 392 -166
rect 392 -167 393 -166
rect 393 -167 394 -166
rect 394 -167 395 -166
rect 395 -167 396 -166
rect 396 -167 397 -166
rect 397 -167 398 -166
rect 398 -167 399 -166
rect 399 -167 400 -166
rect 400 -167 401 -166
rect 401 -167 402 -166
rect 402 -167 403 -166
rect 403 -167 404 -166
rect 404 -167 405 -166
rect 405 -167 406 -166
rect 406 -167 407 -166
rect 407 -167 408 -166
rect 408 -167 409 -166
rect 409 -167 410 -166
rect 410 -167 411 -166
rect 411 -167 412 -166
rect 412 -167 413 -166
rect 413 -167 414 -166
rect 414 -167 415 -166
rect 415 -167 416 -166
rect 416 -167 417 -166
rect 417 -167 418 -166
rect 418 -167 419 -166
rect 419 -167 420 -166
rect 420 -167 421 -166
rect 421 -167 422 -166
rect 422 -167 423 -166
rect 423 -167 424 -166
rect 424 -167 425 -166
rect 425 -167 426 -166
rect 426 -167 427 -166
rect 427 -167 428 -166
rect 428 -167 429 -166
rect 429 -167 430 -166
rect 430 -167 431 -166
rect 431 -167 432 -166
rect 432 -167 433 -166
rect 433 -167 434 -166
rect 434 -167 435 -166
rect 435 -167 436 -166
rect 436 -167 437 -166
rect 437 -167 438 -166
rect 438 -167 439 -166
rect 439 -167 440 -166
rect 440 -167 441 -166
rect 441 -167 442 -166
rect 442 -167 443 -166
rect 443 -167 444 -166
rect 444 -167 445 -166
rect 445 -167 446 -166
rect 446 -167 447 -166
rect 447 -167 448 -166
rect 448 -167 449 -166
rect 449 -167 450 -166
rect 450 -167 451 -166
rect 451 -167 452 -166
rect 452 -167 453 -166
rect 453 -167 454 -166
rect 454 -167 455 -166
rect 455 -167 456 -166
rect 456 -167 457 -166
rect 457 -167 458 -166
rect 458 -167 459 -166
rect 459 -167 460 -166
rect 460 -167 461 -166
rect 461 -167 462 -166
rect 462 -167 463 -166
rect 463 -167 464 -166
rect 464 -167 465 -166
rect 465 -167 466 -166
rect 466 -167 467 -166
rect 467 -167 468 -166
rect 468 -167 469 -166
rect 469 -167 470 -166
rect 470 -167 471 -166
rect 471 -167 472 -166
rect 472 -167 473 -166
rect 473 -167 474 -166
rect 474 -167 475 -166
rect 475 -167 476 -166
rect 476 -167 477 -166
rect 477 -167 478 -166
rect 478 -167 479 -166
rect 479 -167 480 -166
rect 2 -168 3 -167
rect 3 -168 4 -167
rect 4 -168 5 -167
rect 5 -168 6 -167
rect 6 -168 7 -167
rect 7 -168 8 -167
rect 8 -168 9 -167
rect 9 -168 10 -167
rect 10 -168 11 -167
rect 11 -168 12 -167
rect 12 -168 13 -167
rect 13 -168 14 -167
rect 14 -168 15 -167
rect 15 -168 16 -167
rect 16 -168 17 -167
rect 17 -168 18 -167
rect 18 -168 19 -167
rect 19 -168 20 -167
rect 20 -168 21 -167
rect 21 -168 22 -167
rect 22 -168 23 -167
rect 23 -168 24 -167
rect 24 -168 25 -167
rect 25 -168 26 -167
rect 26 -168 27 -167
rect 27 -168 28 -167
rect 28 -168 29 -167
rect 29 -168 30 -167
rect 30 -168 31 -167
rect 31 -168 32 -167
rect 32 -168 33 -167
rect 33 -168 34 -167
rect 34 -168 35 -167
rect 35 -168 36 -167
rect 36 -168 37 -167
rect 37 -168 38 -167
rect 38 -168 39 -167
rect 39 -168 40 -167
rect 40 -168 41 -167
rect 41 -168 42 -167
rect 42 -168 43 -167
rect 43 -168 44 -167
rect 44 -168 45 -167
rect 45 -168 46 -167
rect 46 -168 47 -167
rect 47 -168 48 -167
rect 48 -168 49 -167
rect 49 -168 50 -167
rect 50 -168 51 -167
rect 51 -168 52 -167
rect 52 -168 53 -167
rect 53 -168 54 -167
rect 54 -168 55 -167
rect 55 -168 56 -167
rect 56 -168 57 -167
rect 57 -168 58 -167
rect 58 -168 59 -167
rect 59 -168 60 -167
rect 60 -168 61 -167
rect 61 -168 62 -167
rect 62 -168 63 -167
rect 63 -168 64 -167
rect 64 -168 65 -167
rect 65 -168 66 -167
rect 66 -168 67 -167
rect 67 -168 68 -167
rect 68 -168 69 -167
rect 69 -168 70 -167
rect 70 -168 71 -167
rect 71 -168 72 -167
rect 72 -168 73 -167
rect 73 -168 74 -167
rect 74 -168 75 -167
rect 75 -168 76 -167
rect 76 -168 77 -167
rect 77 -168 78 -167
rect 78 -168 79 -167
rect 79 -168 80 -167
rect 80 -168 81 -167
rect 81 -168 82 -167
rect 82 -168 83 -167
rect 83 -168 84 -167
rect 84 -168 85 -167
rect 85 -168 86 -167
rect 86 -168 87 -167
rect 87 -168 88 -167
rect 88 -168 89 -167
rect 89 -168 90 -167
rect 90 -168 91 -167
rect 91 -168 92 -167
rect 92 -168 93 -167
rect 93 -168 94 -167
rect 94 -168 95 -167
rect 95 -168 96 -167
rect 96 -168 97 -167
rect 97 -168 98 -167
rect 98 -168 99 -167
rect 99 -168 100 -167
rect 100 -168 101 -167
rect 101 -168 102 -167
rect 102 -168 103 -167
rect 103 -168 104 -167
rect 104 -168 105 -167
rect 105 -168 106 -167
rect 106 -168 107 -167
rect 107 -168 108 -167
rect 108 -168 109 -167
rect 109 -168 110 -167
rect 110 -168 111 -167
rect 111 -168 112 -167
rect 112 -168 113 -167
rect 113 -168 114 -167
rect 114 -168 115 -167
rect 115 -168 116 -167
rect 116 -168 117 -167
rect 117 -168 118 -167
rect 118 -168 119 -167
rect 119 -168 120 -167
rect 120 -168 121 -167
rect 121 -168 122 -167
rect 122 -168 123 -167
rect 123 -168 124 -167
rect 124 -168 125 -167
rect 125 -168 126 -167
rect 126 -168 127 -167
rect 127 -168 128 -167
rect 128 -168 129 -167
rect 129 -168 130 -167
rect 130 -168 131 -167
rect 131 -168 132 -167
rect 132 -168 133 -167
rect 133 -168 134 -167
rect 134 -168 135 -167
rect 135 -168 136 -167
rect 136 -168 137 -167
rect 137 -168 138 -167
rect 138 -168 139 -167
rect 139 -168 140 -167
rect 140 -168 141 -167
rect 141 -168 142 -167
rect 142 -168 143 -167
rect 143 -168 144 -167
rect 144 -168 145 -167
rect 145 -168 146 -167
rect 146 -168 147 -167
rect 147 -168 148 -167
rect 148 -168 149 -167
rect 149 -168 150 -167
rect 150 -168 151 -167
rect 151 -168 152 -167
rect 152 -168 153 -167
rect 153 -168 154 -167
rect 154 -168 155 -167
rect 155 -168 156 -167
rect 156 -168 157 -167
rect 157 -168 158 -167
rect 158 -168 159 -167
rect 159 -168 160 -167
rect 160 -168 161 -167
rect 161 -168 162 -167
rect 162 -168 163 -167
rect 163 -168 164 -167
rect 164 -168 165 -167
rect 165 -168 166 -167
rect 166 -168 167 -167
rect 167 -168 168 -167
rect 168 -168 169 -167
rect 169 -168 170 -167
rect 170 -168 171 -167
rect 171 -168 172 -167
rect 172 -168 173 -167
rect 173 -168 174 -167
rect 174 -168 175 -167
rect 175 -168 176 -167
rect 176 -168 177 -167
rect 177 -168 178 -167
rect 178 -168 179 -167
rect 179 -168 180 -167
rect 180 -168 181 -167
rect 181 -168 182 -167
rect 182 -168 183 -167
rect 183 -168 184 -167
rect 184 -168 185 -167
rect 185 -168 186 -167
rect 186 -168 187 -167
rect 187 -168 188 -167
rect 188 -168 189 -167
rect 189 -168 190 -167
rect 190 -168 191 -167
rect 191 -168 192 -167
rect 192 -168 193 -167
rect 193 -168 194 -167
rect 194 -168 195 -167
rect 195 -168 196 -167
rect 196 -168 197 -167
rect 197 -168 198 -167
rect 198 -168 199 -167
rect 199 -168 200 -167
rect 200 -168 201 -167
rect 201 -168 202 -167
rect 202 -168 203 -167
rect 203 -168 204 -167
rect 204 -168 205 -167
rect 205 -168 206 -167
rect 206 -168 207 -167
rect 207 -168 208 -167
rect 208 -168 209 -167
rect 209 -168 210 -167
rect 210 -168 211 -167
rect 211 -168 212 -167
rect 212 -168 213 -167
rect 213 -168 214 -167
rect 214 -168 215 -167
rect 215 -168 216 -167
rect 216 -168 217 -167
rect 217 -168 218 -167
rect 218 -168 219 -167
rect 219 -168 220 -167
rect 220 -168 221 -167
rect 221 -168 222 -167
rect 222 -168 223 -167
rect 223 -168 224 -167
rect 224 -168 225 -167
rect 225 -168 226 -167
rect 226 -168 227 -167
rect 227 -168 228 -167
rect 228 -168 229 -167
rect 229 -168 230 -167
rect 230 -168 231 -167
rect 231 -168 232 -167
rect 232 -168 233 -167
rect 233 -168 234 -167
rect 234 -168 235 -167
rect 235 -168 236 -167
rect 236 -168 237 -167
rect 237 -168 238 -167
rect 238 -168 239 -167
rect 239 -168 240 -167
rect 240 -168 241 -167
rect 241 -168 242 -167
rect 242 -168 243 -167
rect 243 -168 244 -167
rect 244 -168 245 -167
rect 245 -168 246 -167
rect 246 -168 247 -167
rect 247 -168 248 -167
rect 248 -168 249 -167
rect 249 -168 250 -167
rect 250 -168 251 -167
rect 251 -168 252 -167
rect 252 -168 253 -167
rect 253 -168 254 -167
rect 254 -168 255 -167
rect 255 -168 256 -167
rect 256 -168 257 -167
rect 257 -168 258 -167
rect 258 -168 259 -167
rect 259 -168 260 -167
rect 260 -168 261 -167
rect 261 -168 262 -167
rect 262 -168 263 -167
rect 263 -168 264 -167
rect 264 -168 265 -167
rect 265 -168 266 -167
rect 266 -168 267 -167
rect 267 -168 268 -167
rect 268 -168 269 -167
rect 269 -168 270 -167
rect 270 -168 271 -167
rect 271 -168 272 -167
rect 272 -168 273 -167
rect 273 -168 274 -167
rect 274 -168 275 -167
rect 275 -168 276 -167
rect 276 -168 277 -167
rect 277 -168 278 -167
rect 278 -168 279 -167
rect 279 -168 280 -167
rect 280 -168 281 -167
rect 281 -168 282 -167
rect 282 -168 283 -167
rect 283 -168 284 -167
rect 284 -168 285 -167
rect 285 -168 286 -167
rect 286 -168 287 -167
rect 287 -168 288 -167
rect 288 -168 289 -167
rect 289 -168 290 -167
rect 290 -168 291 -167
rect 291 -168 292 -167
rect 292 -168 293 -167
rect 293 -168 294 -167
rect 294 -168 295 -167
rect 295 -168 296 -167
rect 296 -168 297 -167
rect 297 -168 298 -167
rect 298 -168 299 -167
rect 299 -168 300 -167
rect 300 -168 301 -167
rect 301 -168 302 -167
rect 302 -168 303 -167
rect 303 -168 304 -167
rect 304 -168 305 -167
rect 305 -168 306 -167
rect 306 -168 307 -167
rect 307 -168 308 -167
rect 308 -168 309 -167
rect 309 -168 310 -167
rect 310 -168 311 -167
rect 311 -168 312 -167
rect 312 -168 313 -167
rect 313 -168 314 -167
rect 314 -168 315 -167
rect 315 -168 316 -167
rect 316 -168 317 -167
rect 317 -168 318 -167
rect 318 -168 319 -167
rect 319 -168 320 -167
rect 320 -168 321 -167
rect 321 -168 322 -167
rect 322 -168 323 -167
rect 323 -168 324 -167
rect 324 -168 325 -167
rect 325 -168 326 -167
rect 326 -168 327 -167
rect 327 -168 328 -167
rect 328 -168 329 -167
rect 329 -168 330 -167
rect 330 -168 331 -167
rect 331 -168 332 -167
rect 332 -168 333 -167
rect 333 -168 334 -167
rect 334 -168 335 -167
rect 335 -168 336 -167
rect 336 -168 337 -167
rect 337 -168 338 -167
rect 338 -168 339 -167
rect 339 -168 340 -167
rect 340 -168 341 -167
rect 341 -168 342 -167
rect 342 -168 343 -167
rect 343 -168 344 -167
rect 344 -168 345 -167
rect 345 -168 346 -167
rect 346 -168 347 -167
rect 347 -168 348 -167
rect 348 -168 349 -167
rect 349 -168 350 -167
rect 350 -168 351 -167
rect 351 -168 352 -167
rect 352 -168 353 -167
rect 353 -168 354 -167
rect 354 -168 355 -167
rect 355 -168 356 -167
rect 356 -168 357 -167
rect 357 -168 358 -167
rect 358 -168 359 -167
rect 359 -168 360 -167
rect 360 -168 361 -167
rect 361 -168 362 -167
rect 362 -168 363 -167
rect 363 -168 364 -167
rect 364 -168 365 -167
rect 365 -168 366 -167
rect 366 -168 367 -167
rect 367 -168 368 -167
rect 368 -168 369 -167
rect 369 -168 370 -167
rect 370 -168 371 -167
rect 371 -168 372 -167
rect 372 -168 373 -167
rect 373 -168 374 -167
rect 374 -168 375 -167
rect 375 -168 376 -167
rect 376 -168 377 -167
rect 377 -168 378 -167
rect 378 -168 379 -167
rect 379 -168 380 -167
rect 380 -168 381 -167
rect 381 -168 382 -167
rect 382 -168 383 -167
rect 383 -168 384 -167
rect 384 -168 385 -167
rect 385 -168 386 -167
rect 386 -168 387 -167
rect 387 -168 388 -167
rect 388 -168 389 -167
rect 389 -168 390 -167
rect 390 -168 391 -167
rect 391 -168 392 -167
rect 392 -168 393 -167
rect 393 -168 394 -167
rect 394 -168 395 -167
rect 395 -168 396 -167
rect 396 -168 397 -167
rect 397 -168 398 -167
rect 398 -168 399 -167
rect 399 -168 400 -167
rect 400 -168 401 -167
rect 401 -168 402 -167
rect 402 -168 403 -167
rect 403 -168 404 -167
rect 404 -168 405 -167
rect 405 -168 406 -167
rect 406 -168 407 -167
rect 407 -168 408 -167
rect 408 -168 409 -167
rect 409 -168 410 -167
rect 410 -168 411 -167
rect 411 -168 412 -167
rect 412 -168 413 -167
rect 413 -168 414 -167
rect 414 -168 415 -167
rect 415 -168 416 -167
rect 416 -168 417 -167
rect 417 -168 418 -167
rect 418 -168 419 -167
rect 419 -168 420 -167
rect 420 -168 421 -167
rect 421 -168 422 -167
rect 422 -168 423 -167
rect 423 -168 424 -167
rect 424 -168 425 -167
rect 425 -168 426 -167
rect 426 -168 427 -167
rect 427 -168 428 -167
rect 428 -168 429 -167
rect 429 -168 430 -167
rect 430 -168 431 -167
rect 431 -168 432 -167
rect 432 -168 433 -167
rect 433 -168 434 -167
rect 434 -168 435 -167
rect 435 -168 436 -167
rect 436 -168 437 -167
rect 437 -168 438 -167
rect 438 -168 439 -167
rect 439 -168 440 -167
rect 440 -168 441 -167
rect 441 -168 442 -167
rect 442 -168 443 -167
rect 443 -168 444 -167
rect 444 -168 445 -167
rect 445 -168 446 -167
rect 446 -168 447 -167
rect 447 -168 448 -167
rect 448 -168 449 -167
rect 449 -168 450 -167
rect 450 -168 451 -167
rect 451 -168 452 -167
rect 452 -168 453 -167
rect 453 -168 454 -167
rect 454 -168 455 -167
rect 455 -168 456 -167
rect 456 -168 457 -167
rect 457 -168 458 -167
rect 458 -168 459 -167
rect 459 -168 460 -167
rect 460 -168 461 -167
rect 461 -168 462 -167
rect 462 -168 463 -167
rect 463 -168 464 -167
rect 464 -168 465 -167
rect 465 -168 466 -167
rect 466 -168 467 -167
rect 467 -168 468 -167
rect 468 -168 469 -167
rect 469 -168 470 -167
rect 470 -168 471 -167
rect 471 -168 472 -167
rect 472 -168 473 -167
rect 473 -168 474 -167
rect 474 -168 475 -167
rect 475 -168 476 -167
rect 476 -168 477 -167
rect 477 -168 478 -167
rect 478 -168 479 -167
rect 479 -168 480 -167
rect 2 -169 3 -168
rect 3 -169 4 -168
rect 4 -169 5 -168
rect 5 -169 6 -168
rect 6 -169 7 -168
rect 7 -169 8 -168
rect 8 -169 9 -168
rect 9 -169 10 -168
rect 10 -169 11 -168
rect 11 -169 12 -168
rect 12 -169 13 -168
rect 13 -169 14 -168
rect 14 -169 15 -168
rect 15 -169 16 -168
rect 16 -169 17 -168
rect 17 -169 18 -168
rect 18 -169 19 -168
rect 19 -169 20 -168
rect 20 -169 21 -168
rect 21 -169 22 -168
rect 22 -169 23 -168
rect 23 -169 24 -168
rect 24 -169 25 -168
rect 25 -169 26 -168
rect 26 -169 27 -168
rect 27 -169 28 -168
rect 28 -169 29 -168
rect 29 -169 30 -168
rect 30 -169 31 -168
rect 31 -169 32 -168
rect 32 -169 33 -168
rect 33 -169 34 -168
rect 34 -169 35 -168
rect 35 -169 36 -168
rect 36 -169 37 -168
rect 37 -169 38 -168
rect 38 -169 39 -168
rect 39 -169 40 -168
rect 40 -169 41 -168
rect 41 -169 42 -168
rect 42 -169 43 -168
rect 43 -169 44 -168
rect 44 -169 45 -168
rect 45 -169 46 -168
rect 46 -169 47 -168
rect 47 -169 48 -168
rect 48 -169 49 -168
rect 49 -169 50 -168
rect 50 -169 51 -168
rect 51 -169 52 -168
rect 52 -169 53 -168
rect 53 -169 54 -168
rect 54 -169 55 -168
rect 55 -169 56 -168
rect 56 -169 57 -168
rect 57 -169 58 -168
rect 58 -169 59 -168
rect 59 -169 60 -168
rect 60 -169 61 -168
rect 61 -169 62 -168
rect 62 -169 63 -168
rect 63 -169 64 -168
rect 64 -169 65 -168
rect 65 -169 66 -168
rect 66 -169 67 -168
rect 67 -169 68 -168
rect 68 -169 69 -168
rect 69 -169 70 -168
rect 70 -169 71 -168
rect 71 -169 72 -168
rect 72 -169 73 -168
rect 73 -169 74 -168
rect 74 -169 75 -168
rect 75 -169 76 -168
rect 76 -169 77 -168
rect 77 -169 78 -168
rect 78 -169 79 -168
rect 79 -169 80 -168
rect 80 -169 81 -168
rect 81 -169 82 -168
rect 82 -169 83 -168
rect 83 -169 84 -168
rect 84 -169 85 -168
rect 85 -169 86 -168
rect 86 -169 87 -168
rect 87 -169 88 -168
rect 88 -169 89 -168
rect 89 -169 90 -168
rect 90 -169 91 -168
rect 91 -169 92 -168
rect 92 -169 93 -168
rect 93 -169 94 -168
rect 94 -169 95 -168
rect 95 -169 96 -168
rect 96 -169 97 -168
rect 97 -169 98 -168
rect 98 -169 99 -168
rect 99 -169 100 -168
rect 100 -169 101 -168
rect 101 -169 102 -168
rect 102 -169 103 -168
rect 103 -169 104 -168
rect 104 -169 105 -168
rect 105 -169 106 -168
rect 106 -169 107 -168
rect 107 -169 108 -168
rect 108 -169 109 -168
rect 109 -169 110 -168
rect 110 -169 111 -168
rect 111 -169 112 -168
rect 112 -169 113 -168
rect 113 -169 114 -168
rect 114 -169 115 -168
rect 115 -169 116 -168
rect 116 -169 117 -168
rect 117 -169 118 -168
rect 118 -169 119 -168
rect 119 -169 120 -168
rect 120 -169 121 -168
rect 121 -169 122 -168
rect 122 -169 123 -168
rect 123 -169 124 -168
rect 124 -169 125 -168
rect 125 -169 126 -168
rect 126 -169 127 -168
rect 127 -169 128 -168
rect 128 -169 129 -168
rect 129 -169 130 -168
rect 130 -169 131 -168
rect 131 -169 132 -168
rect 132 -169 133 -168
rect 133 -169 134 -168
rect 134 -169 135 -168
rect 135 -169 136 -168
rect 136 -169 137 -168
rect 137 -169 138 -168
rect 138 -169 139 -168
rect 139 -169 140 -168
rect 140 -169 141 -168
rect 141 -169 142 -168
rect 142 -169 143 -168
rect 143 -169 144 -168
rect 144 -169 145 -168
rect 145 -169 146 -168
rect 146 -169 147 -168
rect 147 -169 148 -168
rect 148 -169 149 -168
rect 149 -169 150 -168
rect 150 -169 151 -168
rect 151 -169 152 -168
rect 152 -169 153 -168
rect 153 -169 154 -168
rect 154 -169 155 -168
rect 155 -169 156 -168
rect 156 -169 157 -168
rect 157 -169 158 -168
rect 158 -169 159 -168
rect 159 -169 160 -168
rect 160 -169 161 -168
rect 161 -169 162 -168
rect 162 -169 163 -168
rect 163 -169 164 -168
rect 164 -169 165 -168
rect 165 -169 166 -168
rect 166 -169 167 -168
rect 167 -169 168 -168
rect 168 -169 169 -168
rect 169 -169 170 -168
rect 170 -169 171 -168
rect 171 -169 172 -168
rect 172 -169 173 -168
rect 173 -169 174 -168
rect 174 -169 175 -168
rect 175 -169 176 -168
rect 176 -169 177 -168
rect 177 -169 178 -168
rect 178 -169 179 -168
rect 179 -169 180 -168
rect 180 -169 181 -168
rect 181 -169 182 -168
rect 182 -169 183 -168
rect 183 -169 184 -168
rect 184 -169 185 -168
rect 185 -169 186 -168
rect 186 -169 187 -168
rect 187 -169 188 -168
rect 188 -169 189 -168
rect 189 -169 190 -168
rect 190 -169 191 -168
rect 191 -169 192 -168
rect 192 -169 193 -168
rect 193 -169 194 -168
rect 194 -169 195 -168
rect 195 -169 196 -168
rect 196 -169 197 -168
rect 197 -169 198 -168
rect 198 -169 199 -168
rect 199 -169 200 -168
rect 200 -169 201 -168
rect 201 -169 202 -168
rect 202 -169 203 -168
rect 203 -169 204 -168
rect 204 -169 205 -168
rect 205 -169 206 -168
rect 206 -169 207 -168
rect 207 -169 208 -168
rect 208 -169 209 -168
rect 209 -169 210 -168
rect 210 -169 211 -168
rect 211 -169 212 -168
rect 212 -169 213 -168
rect 213 -169 214 -168
rect 214 -169 215 -168
rect 215 -169 216 -168
rect 216 -169 217 -168
rect 217 -169 218 -168
rect 218 -169 219 -168
rect 219 -169 220 -168
rect 220 -169 221 -168
rect 221 -169 222 -168
rect 222 -169 223 -168
rect 223 -169 224 -168
rect 224 -169 225 -168
rect 225 -169 226 -168
rect 226 -169 227 -168
rect 227 -169 228 -168
rect 228 -169 229 -168
rect 229 -169 230 -168
rect 230 -169 231 -168
rect 231 -169 232 -168
rect 232 -169 233 -168
rect 233 -169 234 -168
rect 234 -169 235 -168
rect 235 -169 236 -168
rect 236 -169 237 -168
rect 237 -169 238 -168
rect 238 -169 239 -168
rect 239 -169 240 -168
rect 240 -169 241 -168
rect 241 -169 242 -168
rect 242 -169 243 -168
rect 243 -169 244 -168
rect 244 -169 245 -168
rect 245 -169 246 -168
rect 246 -169 247 -168
rect 247 -169 248 -168
rect 248 -169 249 -168
rect 249 -169 250 -168
rect 250 -169 251 -168
rect 251 -169 252 -168
rect 252 -169 253 -168
rect 253 -169 254 -168
rect 254 -169 255 -168
rect 255 -169 256 -168
rect 256 -169 257 -168
rect 257 -169 258 -168
rect 258 -169 259 -168
rect 259 -169 260 -168
rect 260 -169 261 -168
rect 261 -169 262 -168
rect 262 -169 263 -168
rect 263 -169 264 -168
rect 264 -169 265 -168
rect 265 -169 266 -168
rect 266 -169 267 -168
rect 267 -169 268 -168
rect 268 -169 269 -168
rect 269 -169 270 -168
rect 270 -169 271 -168
rect 271 -169 272 -168
rect 272 -169 273 -168
rect 273 -169 274 -168
rect 274 -169 275 -168
rect 275 -169 276 -168
rect 276 -169 277 -168
rect 277 -169 278 -168
rect 278 -169 279 -168
rect 279 -169 280 -168
rect 280 -169 281 -168
rect 281 -169 282 -168
rect 282 -169 283 -168
rect 283 -169 284 -168
rect 284 -169 285 -168
rect 285 -169 286 -168
rect 286 -169 287 -168
rect 287 -169 288 -168
rect 288 -169 289 -168
rect 289 -169 290 -168
rect 290 -169 291 -168
rect 291 -169 292 -168
rect 292 -169 293 -168
rect 293 -169 294 -168
rect 294 -169 295 -168
rect 295 -169 296 -168
rect 296 -169 297 -168
rect 297 -169 298 -168
rect 298 -169 299 -168
rect 299 -169 300 -168
rect 300 -169 301 -168
rect 301 -169 302 -168
rect 302 -169 303 -168
rect 303 -169 304 -168
rect 304 -169 305 -168
rect 305 -169 306 -168
rect 306 -169 307 -168
rect 307 -169 308 -168
rect 308 -169 309 -168
rect 309 -169 310 -168
rect 310 -169 311 -168
rect 311 -169 312 -168
rect 312 -169 313 -168
rect 313 -169 314 -168
rect 314 -169 315 -168
rect 315 -169 316 -168
rect 316 -169 317 -168
rect 317 -169 318 -168
rect 318 -169 319 -168
rect 319 -169 320 -168
rect 320 -169 321 -168
rect 321 -169 322 -168
rect 322 -169 323 -168
rect 323 -169 324 -168
rect 324 -169 325 -168
rect 325 -169 326 -168
rect 326 -169 327 -168
rect 327 -169 328 -168
rect 328 -169 329 -168
rect 329 -169 330 -168
rect 330 -169 331 -168
rect 331 -169 332 -168
rect 332 -169 333 -168
rect 333 -169 334 -168
rect 334 -169 335 -168
rect 335 -169 336 -168
rect 336 -169 337 -168
rect 337 -169 338 -168
rect 338 -169 339 -168
rect 339 -169 340 -168
rect 340 -169 341 -168
rect 341 -169 342 -168
rect 342 -169 343 -168
rect 343 -169 344 -168
rect 344 -169 345 -168
rect 345 -169 346 -168
rect 346 -169 347 -168
rect 347 -169 348 -168
rect 348 -169 349 -168
rect 349 -169 350 -168
rect 350 -169 351 -168
rect 351 -169 352 -168
rect 352 -169 353 -168
rect 353 -169 354 -168
rect 354 -169 355 -168
rect 355 -169 356 -168
rect 356 -169 357 -168
rect 357 -169 358 -168
rect 358 -169 359 -168
rect 359 -169 360 -168
rect 360 -169 361 -168
rect 361 -169 362 -168
rect 362 -169 363 -168
rect 363 -169 364 -168
rect 364 -169 365 -168
rect 365 -169 366 -168
rect 366 -169 367 -168
rect 367 -169 368 -168
rect 368 -169 369 -168
rect 369 -169 370 -168
rect 370 -169 371 -168
rect 371 -169 372 -168
rect 372 -169 373 -168
rect 373 -169 374 -168
rect 374 -169 375 -168
rect 375 -169 376 -168
rect 376 -169 377 -168
rect 377 -169 378 -168
rect 378 -169 379 -168
rect 379 -169 380 -168
rect 380 -169 381 -168
rect 381 -169 382 -168
rect 382 -169 383 -168
rect 383 -169 384 -168
rect 384 -169 385 -168
rect 385 -169 386 -168
rect 386 -169 387 -168
rect 387 -169 388 -168
rect 388 -169 389 -168
rect 389 -169 390 -168
rect 390 -169 391 -168
rect 391 -169 392 -168
rect 392 -169 393 -168
rect 393 -169 394 -168
rect 394 -169 395 -168
rect 395 -169 396 -168
rect 396 -169 397 -168
rect 397 -169 398 -168
rect 398 -169 399 -168
rect 399 -169 400 -168
rect 400 -169 401 -168
rect 401 -169 402 -168
rect 402 -169 403 -168
rect 403 -169 404 -168
rect 404 -169 405 -168
rect 405 -169 406 -168
rect 406 -169 407 -168
rect 407 -169 408 -168
rect 408 -169 409 -168
rect 409 -169 410 -168
rect 410 -169 411 -168
rect 411 -169 412 -168
rect 412 -169 413 -168
rect 413 -169 414 -168
rect 414 -169 415 -168
rect 415 -169 416 -168
rect 416 -169 417 -168
rect 417 -169 418 -168
rect 418 -169 419 -168
rect 419 -169 420 -168
rect 420 -169 421 -168
rect 421 -169 422 -168
rect 422 -169 423 -168
rect 423 -169 424 -168
rect 424 -169 425 -168
rect 425 -169 426 -168
rect 426 -169 427 -168
rect 427 -169 428 -168
rect 428 -169 429 -168
rect 429 -169 430 -168
rect 430 -169 431 -168
rect 431 -169 432 -168
rect 432 -169 433 -168
rect 433 -169 434 -168
rect 434 -169 435 -168
rect 435 -169 436 -168
rect 436 -169 437 -168
rect 437 -169 438 -168
rect 438 -169 439 -168
rect 439 -169 440 -168
rect 440 -169 441 -168
rect 441 -169 442 -168
rect 442 -169 443 -168
rect 443 -169 444 -168
rect 444 -169 445 -168
rect 445 -169 446 -168
rect 446 -169 447 -168
rect 447 -169 448 -168
rect 448 -169 449 -168
rect 449 -169 450 -168
rect 450 -169 451 -168
rect 451 -169 452 -168
rect 452 -169 453 -168
rect 453 -169 454 -168
rect 454 -169 455 -168
rect 455 -169 456 -168
rect 456 -169 457 -168
rect 457 -169 458 -168
rect 458 -169 459 -168
rect 459 -169 460 -168
rect 460 -169 461 -168
rect 461 -169 462 -168
rect 462 -169 463 -168
rect 463 -169 464 -168
rect 464 -169 465 -168
rect 465 -169 466 -168
rect 466 -169 467 -168
rect 467 -169 468 -168
rect 468 -169 469 -168
rect 469 -169 470 -168
rect 470 -169 471 -168
rect 471 -169 472 -168
rect 472 -169 473 -168
rect 473 -169 474 -168
rect 474 -169 475 -168
rect 475 -169 476 -168
rect 476 -169 477 -168
rect 477 -169 478 -168
rect 478 -169 479 -168
rect 479 -169 480 -168
rect 2 -170 3 -169
rect 3 -170 4 -169
rect 4 -170 5 -169
rect 5 -170 6 -169
rect 6 -170 7 -169
rect 7 -170 8 -169
rect 8 -170 9 -169
rect 9 -170 10 -169
rect 10 -170 11 -169
rect 11 -170 12 -169
rect 12 -170 13 -169
rect 13 -170 14 -169
rect 14 -170 15 -169
rect 15 -170 16 -169
rect 16 -170 17 -169
rect 17 -170 18 -169
rect 18 -170 19 -169
rect 19 -170 20 -169
rect 20 -170 21 -169
rect 21 -170 22 -169
rect 22 -170 23 -169
rect 23 -170 24 -169
rect 24 -170 25 -169
rect 25 -170 26 -169
rect 26 -170 27 -169
rect 27 -170 28 -169
rect 28 -170 29 -169
rect 29 -170 30 -169
rect 30 -170 31 -169
rect 31 -170 32 -169
rect 32 -170 33 -169
rect 33 -170 34 -169
rect 34 -170 35 -169
rect 35 -170 36 -169
rect 36 -170 37 -169
rect 37 -170 38 -169
rect 38 -170 39 -169
rect 39 -170 40 -169
rect 40 -170 41 -169
rect 41 -170 42 -169
rect 42 -170 43 -169
rect 43 -170 44 -169
rect 44 -170 45 -169
rect 45 -170 46 -169
rect 46 -170 47 -169
rect 47 -170 48 -169
rect 48 -170 49 -169
rect 49 -170 50 -169
rect 50 -170 51 -169
rect 51 -170 52 -169
rect 52 -170 53 -169
rect 53 -170 54 -169
rect 54 -170 55 -169
rect 55 -170 56 -169
rect 56 -170 57 -169
rect 57 -170 58 -169
rect 58 -170 59 -169
rect 59 -170 60 -169
rect 60 -170 61 -169
rect 61 -170 62 -169
rect 62 -170 63 -169
rect 63 -170 64 -169
rect 64 -170 65 -169
rect 65 -170 66 -169
rect 66 -170 67 -169
rect 67 -170 68 -169
rect 68 -170 69 -169
rect 69 -170 70 -169
rect 70 -170 71 -169
rect 71 -170 72 -169
rect 72 -170 73 -169
rect 73 -170 74 -169
rect 74 -170 75 -169
rect 75 -170 76 -169
rect 76 -170 77 -169
rect 77 -170 78 -169
rect 78 -170 79 -169
rect 79 -170 80 -169
rect 80 -170 81 -169
rect 81 -170 82 -169
rect 82 -170 83 -169
rect 83 -170 84 -169
rect 84 -170 85 -169
rect 85 -170 86 -169
rect 86 -170 87 -169
rect 87 -170 88 -169
rect 88 -170 89 -169
rect 89 -170 90 -169
rect 90 -170 91 -169
rect 91 -170 92 -169
rect 92 -170 93 -169
rect 93 -170 94 -169
rect 94 -170 95 -169
rect 95 -170 96 -169
rect 96 -170 97 -169
rect 97 -170 98 -169
rect 98 -170 99 -169
rect 99 -170 100 -169
rect 100 -170 101 -169
rect 101 -170 102 -169
rect 102 -170 103 -169
rect 103 -170 104 -169
rect 104 -170 105 -169
rect 105 -170 106 -169
rect 106 -170 107 -169
rect 107 -170 108 -169
rect 108 -170 109 -169
rect 109 -170 110 -169
rect 110 -170 111 -169
rect 111 -170 112 -169
rect 112 -170 113 -169
rect 113 -170 114 -169
rect 114 -170 115 -169
rect 115 -170 116 -169
rect 116 -170 117 -169
rect 117 -170 118 -169
rect 118 -170 119 -169
rect 119 -170 120 -169
rect 120 -170 121 -169
rect 121 -170 122 -169
rect 122 -170 123 -169
rect 123 -170 124 -169
rect 124 -170 125 -169
rect 125 -170 126 -169
rect 126 -170 127 -169
rect 127 -170 128 -169
rect 128 -170 129 -169
rect 129 -170 130 -169
rect 130 -170 131 -169
rect 131 -170 132 -169
rect 132 -170 133 -169
rect 133 -170 134 -169
rect 134 -170 135 -169
rect 135 -170 136 -169
rect 136 -170 137 -169
rect 137 -170 138 -169
rect 138 -170 139 -169
rect 139 -170 140 -169
rect 140 -170 141 -169
rect 141 -170 142 -169
rect 142 -170 143 -169
rect 143 -170 144 -169
rect 144 -170 145 -169
rect 145 -170 146 -169
rect 146 -170 147 -169
rect 147 -170 148 -169
rect 148 -170 149 -169
rect 149 -170 150 -169
rect 150 -170 151 -169
rect 151 -170 152 -169
rect 152 -170 153 -169
rect 153 -170 154 -169
rect 154 -170 155 -169
rect 155 -170 156 -169
rect 156 -170 157 -169
rect 157 -170 158 -169
rect 158 -170 159 -169
rect 159 -170 160 -169
rect 160 -170 161 -169
rect 161 -170 162 -169
rect 162 -170 163 -169
rect 163 -170 164 -169
rect 164 -170 165 -169
rect 165 -170 166 -169
rect 166 -170 167 -169
rect 167 -170 168 -169
rect 168 -170 169 -169
rect 169 -170 170 -169
rect 170 -170 171 -169
rect 171 -170 172 -169
rect 172 -170 173 -169
rect 173 -170 174 -169
rect 174 -170 175 -169
rect 175 -170 176 -169
rect 176 -170 177 -169
rect 177 -170 178 -169
rect 178 -170 179 -169
rect 179 -170 180 -169
rect 180 -170 181 -169
rect 181 -170 182 -169
rect 182 -170 183 -169
rect 183 -170 184 -169
rect 184 -170 185 -169
rect 185 -170 186 -169
rect 186 -170 187 -169
rect 187 -170 188 -169
rect 188 -170 189 -169
rect 189 -170 190 -169
rect 190 -170 191 -169
rect 191 -170 192 -169
rect 192 -170 193 -169
rect 193 -170 194 -169
rect 194 -170 195 -169
rect 195 -170 196 -169
rect 196 -170 197 -169
rect 197 -170 198 -169
rect 198 -170 199 -169
rect 199 -170 200 -169
rect 200 -170 201 -169
rect 201 -170 202 -169
rect 202 -170 203 -169
rect 203 -170 204 -169
rect 204 -170 205 -169
rect 205 -170 206 -169
rect 206 -170 207 -169
rect 207 -170 208 -169
rect 208 -170 209 -169
rect 209 -170 210 -169
rect 210 -170 211 -169
rect 211 -170 212 -169
rect 212 -170 213 -169
rect 213 -170 214 -169
rect 214 -170 215 -169
rect 215 -170 216 -169
rect 216 -170 217 -169
rect 217 -170 218 -169
rect 218 -170 219 -169
rect 219 -170 220 -169
rect 220 -170 221 -169
rect 221 -170 222 -169
rect 222 -170 223 -169
rect 223 -170 224 -169
rect 224 -170 225 -169
rect 225 -170 226 -169
rect 226 -170 227 -169
rect 227 -170 228 -169
rect 228 -170 229 -169
rect 229 -170 230 -169
rect 230 -170 231 -169
rect 231 -170 232 -169
rect 232 -170 233 -169
rect 233 -170 234 -169
rect 234 -170 235 -169
rect 235 -170 236 -169
rect 236 -170 237 -169
rect 237 -170 238 -169
rect 238 -170 239 -169
rect 239 -170 240 -169
rect 240 -170 241 -169
rect 241 -170 242 -169
rect 242 -170 243 -169
rect 243 -170 244 -169
rect 244 -170 245 -169
rect 245 -170 246 -169
rect 246 -170 247 -169
rect 247 -170 248 -169
rect 248 -170 249 -169
rect 249 -170 250 -169
rect 250 -170 251 -169
rect 251 -170 252 -169
rect 252 -170 253 -169
rect 253 -170 254 -169
rect 254 -170 255 -169
rect 255 -170 256 -169
rect 256 -170 257 -169
rect 257 -170 258 -169
rect 258 -170 259 -169
rect 259 -170 260 -169
rect 260 -170 261 -169
rect 261 -170 262 -169
rect 262 -170 263 -169
rect 263 -170 264 -169
rect 264 -170 265 -169
rect 265 -170 266 -169
rect 266 -170 267 -169
rect 267 -170 268 -169
rect 268 -170 269 -169
rect 269 -170 270 -169
rect 270 -170 271 -169
rect 271 -170 272 -169
rect 272 -170 273 -169
rect 273 -170 274 -169
rect 274 -170 275 -169
rect 275 -170 276 -169
rect 276 -170 277 -169
rect 277 -170 278 -169
rect 278 -170 279 -169
rect 279 -170 280 -169
rect 280 -170 281 -169
rect 281 -170 282 -169
rect 282 -170 283 -169
rect 283 -170 284 -169
rect 284 -170 285 -169
rect 285 -170 286 -169
rect 286 -170 287 -169
rect 287 -170 288 -169
rect 288 -170 289 -169
rect 289 -170 290 -169
rect 290 -170 291 -169
rect 291 -170 292 -169
rect 292 -170 293 -169
rect 293 -170 294 -169
rect 294 -170 295 -169
rect 295 -170 296 -169
rect 296 -170 297 -169
rect 297 -170 298 -169
rect 298 -170 299 -169
rect 299 -170 300 -169
rect 300 -170 301 -169
rect 301 -170 302 -169
rect 302 -170 303 -169
rect 303 -170 304 -169
rect 304 -170 305 -169
rect 305 -170 306 -169
rect 306 -170 307 -169
rect 307 -170 308 -169
rect 308 -170 309 -169
rect 309 -170 310 -169
rect 310 -170 311 -169
rect 311 -170 312 -169
rect 312 -170 313 -169
rect 313 -170 314 -169
rect 314 -170 315 -169
rect 315 -170 316 -169
rect 316 -170 317 -169
rect 317 -170 318 -169
rect 318 -170 319 -169
rect 319 -170 320 -169
rect 320 -170 321 -169
rect 321 -170 322 -169
rect 322 -170 323 -169
rect 323 -170 324 -169
rect 324 -170 325 -169
rect 325 -170 326 -169
rect 326 -170 327 -169
rect 327 -170 328 -169
rect 328 -170 329 -169
rect 329 -170 330 -169
rect 330 -170 331 -169
rect 331 -170 332 -169
rect 332 -170 333 -169
rect 333 -170 334 -169
rect 334 -170 335 -169
rect 335 -170 336 -169
rect 336 -170 337 -169
rect 337 -170 338 -169
rect 338 -170 339 -169
rect 339 -170 340 -169
rect 340 -170 341 -169
rect 341 -170 342 -169
rect 342 -170 343 -169
rect 343 -170 344 -169
rect 344 -170 345 -169
rect 345 -170 346 -169
rect 346 -170 347 -169
rect 347 -170 348 -169
rect 348 -170 349 -169
rect 349 -170 350 -169
rect 350 -170 351 -169
rect 351 -170 352 -169
rect 352 -170 353 -169
rect 353 -170 354 -169
rect 354 -170 355 -169
rect 355 -170 356 -169
rect 356 -170 357 -169
rect 357 -170 358 -169
rect 358 -170 359 -169
rect 359 -170 360 -169
rect 360 -170 361 -169
rect 361 -170 362 -169
rect 362 -170 363 -169
rect 363 -170 364 -169
rect 364 -170 365 -169
rect 365 -170 366 -169
rect 366 -170 367 -169
rect 367 -170 368 -169
rect 368 -170 369 -169
rect 369 -170 370 -169
rect 370 -170 371 -169
rect 371 -170 372 -169
rect 372 -170 373 -169
rect 373 -170 374 -169
rect 374 -170 375 -169
rect 375 -170 376 -169
rect 376 -170 377 -169
rect 377 -170 378 -169
rect 378 -170 379 -169
rect 379 -170 380 -169
rect 380 -170 381 -169
rect 381 -170 382 -169
rect 382 -170 383 -169
rect 383 -170 384 -169
rect 384 -170 385 -169
rect 385 -170 386 -169
rect 386 -170 387 -169
rect 387 -170 388 -169
rect 388 -170 389 -169
rect 389 -170 390 -169
rect 390 -170 391 -169
rect 391 -170 392 -169
rect 392 -170 393 -169
rect 393 -170 394 -169
rect 394 -170 395 -169
rect 395 -170 396 -169
rect 396 -170 397 -169
rect 397 -170 398 -169
rect 398 -170 399 -169
rect 399 -170 400 -169
rect 400 -170 401 -169
rect 401 -170 402 -169
rect 402 -170 403 -169
rect 403 -170 404 -169
rect 404 -170 405 -169
rect 405 -170 406 -169
rect 406 -170 407 -169
rect 407 -170 408 -169
rect 408 -170 409 -169
rect 409 -170 410 -169
rect 410 -170 411 -169
rect 411 -170 412 -169
rect 412 -170 413 -169
rect 413 -170 414 -169
rect 414 -170 415 -169
rect 415 -170 416 -169
rect 416 -170 417 -169
rect 417 -170 418 -169
rect 418 -170 419 -169
rect 419 -170 420 -169
rect 420 -170 421 -169
rect 421 -170 422 -169
rect 422 -170 423 -169
rect 423 -170 424 -169
rect 424 -170 425 -169
rect 425 -170 426 -169
rect 426 -170 427 -169
rect 427 -170 428 -169
rect 428 -170 429 -169
rect 429 -170 430 -169
rect 430 -170 431 -169
rect 431 -170 432 -169
rect 432 -170 433 -169
rect 433 -170 434 -169
rect 434 -170 435 -169
rect 435 -170 436 -169
rect 436 -170 437 -169
rect 437 -170 438 -169
rect 438 -170 439 -169
rect 439 -170 440 -169
rect 440 -170 441 -169
rect 441 -170 442 -169
rect 442 -170 443 -169
rect 443 -170 444 -169
rect 444 -170 445 -169
rect 445 -170 446 -169
rect 446 -170 447 -169
rect 447 -170 448 -169
rect 448 -170 449 -169
rect 449 -170 450 -169
rect 450 -170 451 -169
rect 451 -170 452 -169
rect 452 -170 453 -169
rect 453 -170 454 -169
rect 454 -170 455 -169
rect 455 -170 456 -169
rect 456 -170 457 -169
rect 457 -170 458 -169
rect 458 -170 459 -169
rect 459 -170 460 -169
rect 460 -170 461 -169
rect 461 -170 462 -169
rect 462 -170 463 -169
rect 463 -170 464 -169
rect 464 -170 465 -169
rect 465 -170 466 -169
rect 466 -170 467 -169
rect 467 -170 468 -169
rect 468 -170 469 -169
rect 469 -170 470 -169
rect 470 -170 471 -169
rect 471 -170 472 -169
rect 472 -170 473 -169
rect 473 -170 474 -169
rect 474 -170 475 -169
rect 475 -170 476 -169
rect 476 -170 477 -169
rect 477 -170 478 -169
rect 478 -170 479 -169
rect 479 -170 480 -169
rect 2 -171 3 -170
rect 3 -171 4 -170
rect 4 -171 5 -170
rect 5 -171 6 -170
rect 6 -171 7 -170
rect 7 -171 8 -170
rect 8 -171 9 -170
rect 9 -171 10 -170
rect 10 -171 11 -170
rect 11 -171 12 -170
rect 12 -171 13 -170
rect 13 -171 14 -170
rect 14 -171 15 -170
rect 15 -171 16 -170
rect 16 -171 17 -170
rect 17 -171 18 -170
rect 18 -171 19 -170
rect 19 -171 20 -170
rect 20 -171 21 -170
rect 21 -171 22 -170
rect 22 -171 23 -170
rect 23 -171 24 -170
rect 24 -171 25 -170
rect 25 -171 26 -170
rect 26 -171 27 -170
rect 27 -171 28 -170
rect 28 -171 29 -170
rect 29 -171 30 -170
rect 30 -171 31 -170
rect 31 -171 32 -170
rect 32 -171 33 -170
rect 33 -171 34 -170
rect 34 -171 35 -170
rect 35 -171 36 -170
rect 36 -171 37 -170
rect 37 -171 38 -170
rect 38 -171 39 -170
rect 39 -171 40 -170
rect 40 -171 41 -170
rect 41 -171 42 -170
rect 42 -171 43 -170
rect 43 -171 44 -170
rect 44 -171 45 -170
rect 45 -171 46 -170
rect 46 -171 47 -170
rect 47 -171 48 -170
rect 48 -171 49 -170
rect 49 -171 50 -170
rect 50 -171 51 -170
rect 51 -171 52 -170
rect 52 -171 53 -170
rect 53 -171 54 -170
rect 54 -171 55 -170
rect 55 -171 56 -170
rect 56 -171 57 -170
rect 57 -171 58 -170
rect 58 -171 59 -170
rect 59 -171 60 -170
rect 60 -171 61 -170
rect 61 -171 62 -170
rect 62 -171 63 -170
rect 63 -171 64 -170
rect 64 -171 65 -170
rect 65 -171 66 -170
rect 66 -171 67 -170
rect 67 -171 68 -170
rect 68 -171 69 -170
rect 69 -171 70 -170
rect 70 -171 71 -170
rect 71 -171 72 -170
rect 72 -171 73 -170
rect 73 -171 74 -170
rect 74 -171 75 -170
rect 75 -171 76 -170
rect 76 -171 77 -170
rect 77 -171 78 -170
rect 78 -171 79 -170
rect 79 -171 80 -170
rect 80 -171 81 -170
rect 81 -171 82 -170
rect 82 -171 83 -170
rect 83 -171 84 -170
rect 84 -171 85 -170
rect 85 -171 86 -170
rect 86 -171 87 -170
rect 87 -171 88 -170
rect 88 -171 89 -170
rect 89 -171 90 -170
rect 90 -171 91 -170
rect 91 -171 92 -170
rect 92 -171 93 -170
rect 93 -171 94 -170
rect 94 -171 95 -170
rect 95 -171 96 -170
rect 96 -171 97 -170
rect 97 -171 98 -170
rect 98 -171 99 -170
rect 99 -171 100 -170
rect 100 -171 101 -170
rect 101 -171 102 -170
rect 102 -171 103 -170
rect 103 -171 104 -170
rect 104 -171 105 -170
rect 105 -171 106 -170
rect 106 -171 107 -170
rect 107 -171 108 -170
rect 108 -171 109 -170
rect 109 -171 110 -170
rect 110 -171 111 -170
rect 111 -171 112 -170
rect 112 -171 113 -170
rect 113 -171 114 -170
rect 114 -171 115 -170
rect 115 -171 116 -170
rect 116 -171 117 -170
rect 117 -171 118 -170
rect 118 -171 119 -170
rect 119 -171 120 -170
rect 120 -171 121 -170
rect 121 -171 122 -170
rect 122 -171 123 -170
rect 123 -171 124 -170
rect 124 -171 125 -170
rect 125 -171 126 -170
rect 126 -171 127 -170
rect 127 -171 128 -170
rect 128 -171 129 -170
rect 129 -171 130 -170
rect 130 -171 131 -170
rect 131 -171 132 -170
rect 132 -171 133 -170
rect 133 -171 134 -170
rect 134 -171 135 -170
rect 135 -171 136 -170
rect 136 -171 137 -170
rect 137 -171 138 -170
rect 138 -171 139 -170
rect 139 -171 140 -170
rect 140 -171 141 -170
rect 141 -171 142 -170
rect 142 -171 143 -170
rect 143 -171 144 -170
rect 144 -171 145 -170
rect 145 -171 146 -170
rect 146 -171 147 -170
rect 147 -171 148 -170
rect 148 -171 149 -170
rect 149 -171 150 -170
rect 150 -171 151 -170
rect 151 -171 152 -170
rect 152 -171 153 -170
rect 153 -171 154 -170
rect 154 -171 155 -170
rect 155 -171 156 -170
rect 156 -171 157 -170
rect 157 -171 158 -170
rect 158 -171 159 -170
rect 159 -171 160 -170
rect 160 -171 161 -170
rect 161 -171 162 -170
rect 162 -171 163 -170
rect 163 -171 164 -170
rect 164 -171 165 -170
rect 165 -171 166 -170
rect 166 -171 167 -170
rect 167 -171 168 -170
rect 168 -171 169 -170
rect 169 -171 170 -170
rect 170 -171 171 -170
rect 171 -171 172 -170
rect 172 -171 173 -170
rect 173 -171 174 -170
rect 174 -171 175 -170
rect 175 -171 176 -170
rect 176 -171 177 -170
rect 177 -171 178 -170
rect 178 -171 179 -170
rect 179 -171 180 -170
rect 180 -171 181 -170
rect 181 -171 182 -170
rect 182 -171 183 -170
rect 183 -171 184 -170
rect 184 -171 185 -170
rect 185 -171 186 -170
rect 186 -171 187 -170
rect 187 -171 188 -170
rect 188 -171 189 -170
rect 189 -171 190 -170
rect 190 -171 191 -170
rect 191 -171 192 -170
rect 192 -171 193 -170
rect 193 -171 194 -170
rect 194 -171 195 -170
rect 195 -171 196 -170
rect 196 -171 197 -170
rect 197 -171 198 -170
rect 198 -171 199 -170
rect 199 -171 200 -170
rect 200 -171 201 -170
rect 201 -171 202 -170
rect 202 -171 203 -170
rect 203 -171 204 -170
rect 204 -171 205 -170
rect 205 -171 206 -170
rect 206 -171 207 -170
rect 207 -171 208 -170
rect 208 -171 209 -170
rect 209 -171 210 -170
rect 210 -171 211 -170
rect 211 -171 212 -170
rect 212 -171 213 -170
rect 213 -171 214 -170
rect 214 -171 215 -170
rect 215 -171 216 -170
rect 216 -171 217 -170
rect 217 -171 218 -170
rect 218 -171 219 -170
rect 219 -171 220 -170
rect 220 -171 221 -170
rect 221 -171 222 -170
rect 222 -171 223 -170
rect 223 -171 224 -170
rect 224 -171 225 -170
rect 225 -171 226 -170
rect 226 -171 227 -170
rect 227 -171 228 -170
rect 228 -171 229 -170
rect 229 -171 230 -170
rect 230 -171 231 -170
rect 231 -171 232 -170
rect 232 -171 233 -170
rect 233 -171 234 -170
rect 234 -171 235 -170
rect 235 -171 236 -170
rect 236 -171 237 -170
rect 237 -171 238 -170
rect 238 -171 239 -170
rect 239 -171 240 -170
rect 240 -171 241 -170
rect 241 -171 242 -170
rect 242 -171 243 -170
rect 243 -171 244 -170
rect 244 -171 245 -170
rect 245 -171 246 -170
rect 246 -171 247 -170
rect 247 -171 248 -170
rect 248 -171 249 -170
rect 249 -171 250 -170
rect 250 -171 251 -170
rect 251 -171 252 -170
rect 252 -171 253 -170
rect 253 -171 254 -170
rect 254 -171 255 -170
rect 255 -171 256 -170
rect 256 -171 257 -170
rect 257 -171 258 -170
rect 258 -171 259 -170
rect 259 -171 260 -170
rect 260 -171 261 -170
rect 261 -171 262 -170
rect 262 -171 263 -170
rect 263 -171 264 -170
rect 264 -171 265 -170
rect 265 -171 266 -170
rect 266 -171 267 -170
rect 267 -171 268 -170
rect 268 -171 269 -170
rect 269 -171 270 -170
rect 270 -171 271 -170
rect 271 -171 272 -170
rect 272 -171 273 -170
rect 273 -171 274 -170
rect 274 -171 275 -170
rect 275 -171 276 -170
rect 276 -171 277 -170
rect 277 -171 278 -170
rect 278 -171 279 -170
rect 279 -171 280 -170
rect 280 -171 281 -170
rect 281 -171 282 -170
rect 282 -171 283 -170
rect 283 -171 284 -170
rect 284 -171 285 -170
rect 285 -171 286 -170
rect 286 -171 287 -170
rect 287 -171 288 -170
rect 288 -171 289 -170
rect 289 -171 290 -170
rect 290 -171 291 -170
rect 291 -171 292 -170
rect 292 -171 293 -170
rect 293 -171 294 -170
rect 294 -171 295 -170
rect 295 -171 296 -170
rect 296 -171 297 -170
rect 297 -171 298 -170
rect 298 -171 299 -170
rect 299 -171 300 -170
rect 300 -171 301 -170
rect 301 -171 302 -170
rect 302 -171 303 -170
rect 303 -171 304 -170
rect 304 -171 305 -170
rect 305 -171 306 -170
rect 306 -171 307 -170
rect 307 -171 308 -170
rect 308 -171 309 -170
rect 309 -171 310 -170
rect 310 -171 311 -170
rect 311 -171 312 -170
rect 312 -171 313 -170
rect 313 -171 314 -170
rect 314 -171 315 -170
rect 315 -171 316 -170
rect 316 -171 317 -170
rect 317 -171 318 -170
rect 318 -171 319 -170
rect 319 -171 320 -170
rect 320 -171 321 -170
rect 321 -171 322 -170
rect 322 -171 323 -170
rect 323 -171 324 -170
rect 324 -171 325 -170
rect 325 -171 326 -170
rect 326 -171 327 -170
rect 327 -171 328 -170
rect 328 -171 329 -170
rect 329 -171 330 -170
rect 330 -171 331 -170
rect 331 -171 332 -170
rect 332 -171 333 -170
rect 333 -171 334 -170
rect 334 -171 335 -170
rect 335 -171 336 -170
rect 336 -171 337 -170
rect 337 -171 338 -170
rect 338 -171 339 -170
rect 339 -171 340 -170
rect 340 -171 341 -170
rect 341 -171 342 -170
rect 342 -171 343 -170
rect 343 -171 344 -170
rect 344 -171 345 -170
rect 345 -171 346 -170
rect 346 -171 347 -170
rect 347 -171 348 -170
rect 348 -171 349 -170
rect 349 -171 350 -170
rect 350 -171 351 -170
rect 351 -171 352 -170
rect 352 -171 353 -170
rect 353 -171 354 -170
rect 354 -171 355 -170
rect 355 -171 356 -170
rect 356 -171 357 -170
rect 357 -171 358 -170
rect 358 -171 359 -170
rect 359 -171 360 -170
rect 360 -171 361 -170
rect 361 -171 362 -170
rect 362 -171 363 -170
rect 363 -171 364 -170
rect 364 -171 365 -170
rect 365 -171 366 -170
rect 366 -171 367 -170
rect 367 -171 368 -170
rect 368 -171 369 -170
rect 369 -171 370 -170
rect 370 -171 371 -170
rect 371 -171 372 -170
rect 372 -171 373 -170
rect 373 -171 374 -170
rect 374 -171 375 -170
rect 375 -171 376 -170
rect 376 -171 377 -170
rect 377 -171 378 -170
rect 378 -171 379 -170
rect 379 -171 380 -170
rect 380 -171 381 -170
rect 381 -171 382 -170
rect 382 -171 383 -170
rect 383 -171 384 -170
rect 384 -171 385 -170
rect 385 -171 386 -170
rect 386 -171 387 -170
rect 387 -171 388 -170
rect 388 -171 389 -170
rect 389 -171 390 -170
rect 390 -171 391 -170
rect 391 -171 392 -170
rect 392 -171 393 -170
rect 393 -171 394 -170
rect 394 -171 395 -170
rect 395 -171 396 -170
rect 396 -171 397 -170
rect 397 -171 398 -170
rect 398 -171 399 -170
rect 399 -171 400 -170
rect 400 -171 401 -170
rect 401 -171 402 -170
rect 402 -171 403 -170
rect 403 -171 404 -170
rect 404 -171 405 -170
rect 405 -171 406 -170
rect 406 -171 407 -170
rect 407 -171 408 -170
rect 408 -171 409 -170
rect 409 -171 410 -170
rect 410 -171 411 -170
rect 411 -171 412 -170
rect 412 -171 413 -170
rect 413 -171 414 -170
rect 414 -171 415 -170
rect 415 -171 416 -170
rect 416 -171 417 -170
rect 417 -171 418 -170
rect 418 -171 419 -170
rect 419 -171 420 -170
rect 420 -171 421 -170
rect 421 -171 422 -170
rect 422 -171 423 -170
rect 423 -171 424 -170
rect 424 -171 425 -170
rect 425 -171 426 -170
rect 426 -171 427 -170
rect 427 -171 428 -170
rect 428 -171 429 -170
rect 429 -171 430 -170
rect 430 -171 431 -170
rect 431 -171 432 -170
rect 432 -171 433 -170
rect 433 -171 434 -170
rect 434 -171 435 -170
rect 435 -171 436 -170
rect 436 -171 437 -170
rect 437 -171 438 -170
rect 438 -171 439 -170
rect 439 -171 440 -170
rect 440 -171 441 -170
rect 441 -171 442 -170
rect 442 -171 443 -170
rect 443 -171 444 -170
rect 444 -171 445 -170
rect 445 -171 446 -170
rect 446 -171 447 -170
rect 447 -171 448 -170
rect 448 -171 449 -170
rect 449 -171 450 -170
rect 450 -171 451 -170
rect 451 -171 452 -170
rect 452 -171 453 -170
rect 453 -171 454 -170
rect 454 -171 455 -170
rect 455 -171 456 -170
rect 456 -171 457 -170
rect 457 -171 458 -170
rect 458 -171 459 -170
rect 459 -171 460 -170
rect 460 -171 461 -170
rect 461 -171 462 -170
rect 462 -171 463 -170
rect 463 -171 464 -170
rect 464 -171 465 -170
rect 465 -171 466 -170
rect 466 -171 467 -170
rect 467 -171 468 -170
rect 468 -171 469 -170
rect 469 -171 470 -170
rect 470 -171 471 -170
rect 471 -171 472 -170
rect 472 -171 473 -170
rect 473 -171 474 -170
rect 474 -171 475 -170
rect 475 -171 476 -170
rect 476 -171 477 -170
rect 477 -171 478 -170
rect 478 -171 479 -170
rect 479 -171 480 -170
rect 2 -172 3 -171
rect 3 -172 4 -171
rect 4 -172 5 -171
rect 5 -172 6 -171
rect 6 -172 7 -171
rect 7 -172 8 -171
rect 8 -172 9 -171
rect 9 -172 10 -171
rect 10 -172 11 -171
rect 11 -172 12 -171
rect 12 -172 13 -171
rect 13 -172 14 -171
rect 14 -172 15 -171
rect 15 -172 16 -171
rect 16 -172 17 -171
rect 17 -172 18 -171
rect 18 -172 19 -171
rect 19 -172 20 -171
rect 20 -172 21 -171
rect 21 -172 22 -171
rect 22 -172 23 -171
rect 23 -172 24 -171
rect 24 -172 25 -171
rect 25 -172 26 -171
rect 26 -172 27 -171
rect 27 -172 28 -171
rect 28 -172 29 -171
rect 29 -172 30 -171
rect 30 -172 31 -171
rect 31 -172 32 -171
rect 32 -172 33 -171
rect 33 -172 34 -171
rect 34 -172 35 -171
rect 35 -172 36 -171
rect 36 -172 37 -171
rect 37 -172 38 -171
rect 38 -172 39 -171
rect 39 -172 40 -171
rect 40 -172 41 -171
rect 41 -172 42 -171
rect 42 -172 43 -171
rect 43 -172 44 -171
rect 44 -172 45 -171
rect 45 -172 46 -171
rect 46 -172 47 -171
rect 47 -172 48 -171
rect 48 -172 49 -171
rect 49 -172 50 -171
rect 50 -172 51 -171
rect 51 -172 52 -171
rect 52 -172 53 -171
rect 53 -172 54 -171
rect 54 -172 55 -171
rect 55 -172 56 -171
rect 56 -172 57 -171
rect 57 -172 58 -171
rect 58 -172 59 -171
rect 59 -172 60 -171
rect 60 -172 61 -171
rect 61 -172 62 -171
rect 62 -172 63 -171
rect 63 -172 64 -171
rect 64 -172 65 -171
rect 65 -172 66 -171
rect 66 -172 67 -171
rect 67 -172 68 -171
rect 68 -172 69 -171
rect 69 -172 70 -171
rect 70 -172 71 -171
rect 71 -172 72 -171
rect 72 -172 73 -171
rect 73 -172 74 -171
rect 74 -172 75 -171
rect 75 -172 76 -171
rect 76 -172 77 -171
rect 77 -172 78 -171
rect 78 -172 79 -171
rect 79 -172 80 -171
rect 80 -172 81 -171
rect 81 -172 82 -171
rect 82 -172 83 -171
rect 83 -172 84 -171
rect 84 -172 85 -171
rect 85 -172 86 -171
rect 86 -172 87 -171
rect 87 -172 88 -171
rect 88 -172 89 -171
rect 89 -172 90 -171
rect 90 -172 91 -171
rect 91 -172 92 -171
rect 92 -172 93 -171
rect 93 -172 94 -171
rect 94 -172 95 -171
rect 95 -172 96 -171
rect 96 -172 97 -171
rect 97 -172 98 -171
rect 98 -172 99 -171
rect 99 -172 100 -171
rect 100 -172 101 -171
rect 101 -172 102 -171
rect 102 -172 103 -171
rect 103 -172 104 -171
rect 104 -172 105 -171
rect 105 -172 106 -171
rect 106 -172 107 -171
rect 107 -172 108 -171
rect 108 -172 109 -171
rect 109 -172 110 -171
rect 110 -172 111 -171
rect 111 -172 112 -171
rect 112 -172 113 -171
rect 113 -172 114 -171
rect 114 -172 115 -171
rect 115 -172 116 -171
rect 116 -172 117 -171
rect 117 -172 118 -171
rect 118 -172 119 -171
rect 119 -172 120 -171
rect 120 -172 121 -171
rect 121 -172 122 -171
rect 122 -172 123 -171
rect 123 -172 124 -171
rect 124 -172 125 -171
rect 125 -172 126 -171
rect 126 -172 127 -171
rect 127 -172 128 -171
rect 128 -172 129 -171
rect 129 -172 130 -171
rect 130 -172 131 -171
rect 131 -172 132 -171
rect 132 -172 133 -171
rect 133 -172 134 -171
rect 134 -172 135 -171
rect 135 -172 136 -171
rect 136 -172 137 -171
rect 137 -172 138 -171
rect 138 -172 139 -171
rect 139 -172 140 -171
rect 140 -172 141 -171
rect 141 -172 142 -171
rect 142 -172 143 -171
rect 143 -172 144 -171
rect 144 -172 145 -171
rect 145 -172 146 -171
rect 146 -172 147 -171
rect 147 -172 148 -171
rect 148 -172 149 -171
rect 149 -172 150 -171
rect 150 -172 151 -171
rect 151 -172 152 -171
rect 152 -172 153 -171
rect 153 -172 154 -171
rect 154 -172 155 -171
rect 155 -172 156 -171
rect 156 -172 157 -171
rect 157 -172 158 -171
rect 158 -172 159 -171
rect 159 -172 160 -171
rect 160 -172 161 -171
rect 161 -172 162 -171
rect 162 -172 163 -171
rect 163 -172 164 -171
rect 164 -172 165 -171
rect 165 -172 166 -171
rect 166 -172 167 -171
rect 167 -172 168 -171
rect 168 -172 169 -171
rect 169 -172 170 -171
rect 170 -172 171 -171
rect 171 -172 172 -171
rect 172 -172 173 -171
rect 173 -172 174 -171
rect 174 -172 175 -171
rect 175 -172 176 -171
rect 176 -172 177 -171
rect 177 -172 178 -171
rect 178 -172 179 -171
rect 179 -172 180 -171
rect 180 -172 181 -171
rect 181 -172 182 -171
rect 182 -172 183 -171
rect 183 -172 184 -171
rect 184 -172 185 -171
rect 185 -172 186 -171
rect 186 -172 187 -171
rect 187 -172 188 -171
rect 188 -172 189 -171
rect 189 -172 190 -171
rect 190 -172 191 -171
rect 191 -172 192 -171
rect 192 -172 193 -171
rect 193 -172 194 -171
rect 194 -172 195 -171
rect 195 -172 196 -171
rect 196 -172 197 -171
rect 197 -172 198 -171
rect 198 -172 199 -171
rect 199 -172 200 -171
rect 200 -172 201 -171
rect 201 -172 202 -171
rect 202 -172 203 -171
rect 203 -172 204 -171
rect 204 -172 205 -171
rect 205 -172 206 -171
rect 206 -172 207 -171
rect 207 -172 208 -171
rect 208 -172 209 -171
rect 209 -172 210 -171
rect 210 -172 211 -171
rect 211 -172 212 -171
rect 212 -172 213 -171
rect 213 -172 214 -171
rect 214 -172 215 -171
rect 215 -172 216 -171
rect 216 -172 217 -171
rect 217 -172 218 -171
rect 218 -172 219 -171
rect 219 -172 220 -171
rect 220 -172 221 -171
rect 221 -172 222 -171
rect 222 -172 223 -171
rect 223 -172 224 -171
rect 224 -172 225 -171
rect 225 -172 226 -171
rect 226 -172 227 -171
rect 227 -172 228 -171
rect 228 -172 229 -171
rect 229 -172 230 -171
rect 230 -172 231 -171
rect 231 -172 232 -171
rect 232 -172 233 -171
rect 233 -172 234 -171
rect 234 -172 235 -171
rect 235 -172 236 -171
rect 236 -172 237 -171
rect 237 -172 238 -171
rect 238 -172 239 -171
rect 239 -172 240 -171
rect 240 -172 241 -171
rect 241 -172 242 -171
rect 242 -172 243 -171
rect 243 -172 244 -171
rect 244 -172 245 -171
rect 245 -172 246 -171
rect 246 -172 247 -171
rect 247 -172 248 -171
rect 248 -172 249 -171
rect 249 -172 250 -171
rect 250 -172 251 -171
rect 251 -172 252 -171
rect 252 -172 253 -171
rect 253 -172 254 -171
rect 254 -172 255 -171
rect 255 -172 256 -171
rect 256 -172 257 -171
rect 257 -172 258 -171
rect 258 -172 259 -171
rect 259 -172 260 -171
rect 260 -172 261 -171
rect 261 -172 262 -171
rect 262 -172 263 -171
rect 263 -172 264 -171
rect 264 -172 265 -171
rect 265 -172 266 -171
rect 266 -172 267 -171
rect 267 -172 268 -171
rect 268 -172 269 -171
rect 269 -172 270 -171
rect 270 -172 271 -171
rect 271 -172 272 -171
rect 272 -172 273 -171
rect 273 -172 274 -171
rect 274 -172 275 -171
rect 275 -172 276 -171
rect 276 -172 277 -171
rect 277 -172 278 -171
rect 278 -172 279 -171
rect 279 -172 280 -171
rect 280 -172 281 -171
rect 281 -172 282 -171
rect 282 -172 283 -171
rect 283 -172 284 -171
rect 284 -172 285 -171
rect 285 -172 286 -171
rect 286 -172 287 -171
rect 287 -172 288 -171
rect 288 -172 289 -171
rect 289 -172 290 -171
rect 290 -172 291 -171
rect 291 -172 292 -171
rect 292 -172 293 -171
rect 293 -172 294 -171
rect 294 -172 295 -171
rect 295 -172 296 -171
rect 296 -172 297 -171
rect 297 -172 298 -171
rect 298 -172 299 -171
rect 299 -172 300 -171
rect 300 -172 301 -171
rect 301 -172 302 -171
rect 302 -172 303 -171
rect 303 -172 304 -171
rect 304 -172 305 -171
rect 305 -172 306 -171
rect 306 -172 307 -171
rect 307 -172 308 -171
rect 308 -172 309 -171
rect 309 -172 310 -171
rect 310 -172 311 -171
rect 311 -172 312 -171
rect 312 -172 313 -171
rect 313 -172 314 -171
rect 314 -172 315 -171
rect 315 -172 316 -171
rect 316 -172 317 -171
rect 317 -172 318 -171
rect 318 -172 319 -171
rect 319 -172 320 -171
rect 320 -172 321 -171
rect 321 -172 322 -171
rect 322 -172 323 -171
rect 323 -172 324 -171
rect 324 -172 325 -171
rect 325 -172 326 -171
rect 326 -172 327 -171
rect 327 -172 328 -171
rect 328 -172 329 -171
rect 329 -172 330 -171
rect 330 -172 331 -171
rect 331 -172 332 -171
rect 332 -172 333 -171
rect 333 -172 334 -171
rect 334 -172 335 -171
rect 335 -172 336 -171
rect 336 -172 337 -171
rect 337 -172 338 -171
rect 338 -172 339 -171
rect 339 -172 340 -171
rect 340 -172 341 -171
rect 341 -172 342 -171
rect 342 -172 343 -171
rect 343 -172 344 -171
rect 344 -172 345 -171
rect 345 -172 346 -171
rect 346 -172 347 -171
rect 347 -172 348 -171
rect 348 -172 349 -171
rect 349 -172 350 -171
rect 350 -172 351 -171
rect 351 -172 352 -171
rect 352 -172 353 -171
rect 353 -172 354 -171
rect 354 -172 355 -171
rect 355 -172 356 -171
rect 356 -172 357 -171
rect 357 -172 358 -171
rect 358 -172 359 -171
rect 359 -172 360 -171
rect 360 -172 361 -171
rect 361 -172 362 -171
rect 362 -172 363 -171
rect 363 -172 364 -171
rect 364 -172 365 -171
rect 365 -172 366 -171
rect 366 -172 367 -171
rect 367 -172 368 -171
rect 368 -172 369 -171
rect 369 -172 370 -171
rect 370 -172 371 -171
rect 371 -172 372 -171
rect 372 -172 373 -171
rect 373 -172 374 -171
rect 374 -172 375 -171
rect 375 -172 376 -171
rect 376 -172 377 -171
rect 377 -172 378 -171
rect 378 -172 379 -171
rect 379 -172 380 -171
rect 380 -172 381 -171
rect 381 -172 382 -171
rect 382 -172 383 -171
rect 383 -172 384 -171
rect 384 -172 385 -171
rect 385 -172 386 -171
rect 386 -172 387 -171
rect 387 -172 388 -171
rect 388 -172 389 -171
rect 389 -172 390 -171
rect 390 -172 391 -171
rect 391 -172 392 -171
rect 392 -172 393 -171
rect 393 -172 394 -171
rect 394 -172 395 -171
rect 395 -172 396 -171
rect 396 -172 397 -171
rect 397 -172 398 -171
rect 398 -172 399 -171
rect 399 -172 400 -171
rect 400 -172 401 -171
rect 401 -172 402 -171
rect 402 -172 403 -171
rect 403 -172 404 -171
rect 404 -172 405 -171
rect 405 -172 406 -171
rect 406 -172 407 -171
rect 407 -172 408 -171
rect 408 -172 409 -171
rect 409 -172 410 -171
rect 410 -172 411 -171
rect 411 -172 412 -171
rect 412 -172 413 -171
rect 413 -172 414 -171
rect 414 -172 415 -171
rect 415 -172 416 -171
rect 416 -172 417 -171
rect 417 -172 418 -171
rect 418 -172 419 -171
rect 419 -172 420 -171
rect 420 -172 421 -171
rect 421 -172 422 -171
rect 422 -172 423 -171
rect 423 -172 424 -171
rect 424 -172 425 -171
rect 425 -172 426 -171
rect 426 -172 427 -171
rect 427 -172 428 -171
rect 428 -172 429 -171
rect 429 -172 430 -171
rect 430 -172 431 -171
rect 431 -172 432 -171
rect 432 -172 433 -171
rect 433 -172 434 -171
rect 434 -172 435 -171
rect 435 -172 436 -171
rect 436 -172 437 -171
rect 437 -172 438 -171
rect 438 -172 439 -171
rect 439 -172 440 -171
rect 440 -172 441 -171
rect 441 -172 442 -171
rect 442 -172 443 -171
rect 443 -172 444 -171
rect 444 -172 445 -171
rect 445 -172 446 -171
rect 446 -172 447 -171
rect 447 -172 448 -171
rect 448 -172 449 -171
rect 449 -172 450 -171
rect 450 -172 451 -171
rect 451 -172 452 -171
rect 452 -172 453 -171
rect 453 -172 454 -171
rect 454 -172 455 -171
rect 455 -172 456 -171
rect 456 -172 457 -171
rect 457 -172 458 -171
rect 458 -172 459 -171
rect 459 -172 460 -171
rect 460 -172 461 -171
rect 461 -172 462 -171
rect 462 -172 463 -171
rect 463 -172 464 -171
rect 464 -172 465 -171
rect 465 -172 466 -171
rect 466 -172 467 -171
rect 467 -172 468 -171
rect 468 -172 469 -171
rect 469 -172 470 -171
rect 470 -172 471 -171
rect 471 -172 472 -171
rect 472 -172 473 -171
rect 473 -172 474 -171
rect 474 -172 475 -171
rect 475 -172 476 -171
rect 476 -172 477 -171
rect 477 -172 478 -171
rect 478 -172 479 -171
rect 479 -172 480 -171
rect 2 -173 3 -172
rect 3 -173 4 -172
rect 4 -173 5 -172
rect 5 -173 6 -172
rect 6 -173 7 -172
rect 7 -173 8 -172
rect 8 -173 9 -172
rect 9 -173 10 -172
rect 10 -173 11 -172
rect 11 -173 12 -172
rect 12 -173 13 -172
rect 13 -173 14 -172
rect 14 -173 15 -172
rect 15 -173 16 -172
rect 16 -173 17 -172
rect 17 -173 18 -172
rect 18 -173 19 -172
rect 19 -173 20 -172
rect 20 -173 21 -172
rect 21 -173 22 -172
rect 22 -173 23 -172
rect 23 -173 24 -172
rect 24 -173 25 -172
rect 25 -173 26 -172
rect 26 -173 27 -172
rect 27 -173 28 -172
rect 28 -173 29 -172
rect 29 -173 30 -172
rect 30 -173 31 -172
rect 31 -173 32 -172
rect 32 -173 33 -172
rect 33 -173 34 -172
rect 34 -173 35 -172
rect 35 -173 36 -172
rect 36 -173 37 -172
rect 37 -173 38 -172
rect 38 -173 39 -172
rect 39 -173 40 -172
rect 40 -173 41 -172
rect 41 -173 42 -172
rect 42 -173 43 -172
rect 43 -173 44 -172
rect 44 -173 45 -172
rect 45 -173 46 -172
rect 46 -173 47 -172
rect 47 -173 48 -172
rect 48 -173 49 -172
rect 49 -173 50 -172
rect 50 -173 51 -172
rect 51 -173 52 -172
rect 52 -173 53 -172
rect 53 -173 54 -172
rect 54 -173 55 -172
rect 55 -173 56 -172
rect 56 -173 57 -172
rect 57 -173 58 -172
rect 58 -173 59 -172
rect 59 -173 60 -172
rect 60 -173 61 -172
rect 61 -173 62 -172
rect 62 -173 63 -172
rect 63 -173 64 -172
rect 64 -173 65 -172
rect 65 -173 66 -172
rect 66 -173 67 -172
rect 67 -173 68 -172
rect 68 -173 69 -172
rect 69 -173 70 -172
rect 70 -173 71 -172
rect 71 -173 72 -172
rect 72 -173 73 -172
rect 73 -173 74 -172
rect 74 -173 75 -172
rect 75 -173 76 -172
rect 76 -173 77 -172
rect 77 -173 78 -172
rect 78 -173 79 -172
rect 79 -173 80 -172
rect 80 -173 81 -172
rect 81 -173 82 -172
rect 82 -173 83 -172
rect 83 -173 84 -172
rect 84 -173 85 -172
rect 85 -173 86 -172
rect 86 -173 87 -172
rect 87 -173 88 -172
rect 88 -173 89 -172
rect 89 -173 90 -172
rect 90 -173 91 -172
rect 91 -173 92 -172
rect 92 -173 93 -172
rect 93 -173 94 -172
rect 94 -173 95 -172
rect 95 -173 96 -172
rect 96 -173 97 -172
rect 97 -173 98 -172
rect 98 -173 99 -172
rect 99 -173 100 -172
rect 100 -173 101 -172
rect 101 -173 102 -172
rect 102 -173 103 -172
rect 103 -173 104 -172
rect 104 -173 105 -172
rect 105 -173 106 -172
rect 106 -173 107 -172
rect 107 -173 108 -172
rect 108 -173 109 -172
rect 109 -173 110 -172
rect 110 -173 111 -172
rect 111 -173 112 -172
rect 112 -173 113 -172
rect 113 -173 114 -172
rect 114 -173 115 -172
rect 115 -173 116 -172
rect 116 -173 117 -172
rect 117 -173 118 -172
rect 118 -173 119 -172
rect 119 -173 120 -172
rect 120 -173 121 -172
rect 121 -173 122 -172
rect 122 -173 123 -172
rect 123 -173 124 -172
rect 124 -173 125 -172
rect 125 -173 126 -172
rect 126 -173 127 -172
rect 127 -173 128 -172
rect 128 -173 129 -172
rect 129 -173 130 -172
rect 130 -173 131 -172
rect 131 -173 132 -172
rect 132 -173 133 -172
rect 133 -173 134 -172
rect 134 -173 135 -172
rect 135 -173 136 -172
rect 136 -173 137 -172
rect 137 -173 138 -172
rect 138 -173 139 -172
rect 139 -173 140 -172
rect 140 -173 141 -172
rect 141 -173 142 -172
rect 142 -173 143 -172
rect 143 -173 144 -172
rect 144 -173 145 -172
rect 145 -173 146 -172
rect 146 -173 147 -172
rect 147 -173 148 -172
rect 148 -173 149 -172
rect 149 -173 150 -172
rect 150 -173 151 -172
rect 151 -173 152 -172
rect 152 -173 153 -172
rect 153 -173 154 -172
rect 154 -173 155 -172
rect 155 -173 156 -172
rect 156 -173 157 -172
rect 157 -173 158 -172
rect 158 -173 159 -172
rect 159 -173 160 -172
rect 160 -173 161 -172
rect 161 -173 162 -172
rect 162 -173 163 -172
rect 163 -173 164 -172
rect 164 -173 165 -172
rect 165 -173 166 -172
rect 166 -173 167 -172
rect 167 -173 168 -172
rect 168 -173 169 -172
rect 169 -173 170 -172
rect 170 -173 171 -172
rect 171 -173 172 -172
rect 172 -173 173 -172
rect 173 -173 174 -172
rect 174 -173 175 -172
rect 175 -173 176 -172
rect 176 -173 177 -172
rect 177 -173 178 -172
rect 178 -173 179 -172
rect 179 -173 180 -172
rect 180 -173 181 -172
rect 181 -173 182 -172
rect 182 -173 183 -172
rect 183 -173 184 -172
rect 184 -173 185 -172
rect 185 -173 186 -172
rect 186 -173 187 -172
rect 187 -173 188 -172
rect 188 -173 189 -172
rect 189 -173 190 -172
rect 190 -173 191 -172
rect 191 -173 192 -172
rect 192 -173 193 -172
rect 193 -173 194 -172
rect 194 -173 195 -172
rect 195 -173 196 -172
rect 196 -173 197 -172
rect 197 -173 198 -172
rect 198 -173 199 -172
rect 199 -173 200 -172
rect 200 -173 201 -172
rect 201 -173 202 -172
rect 202 -173 203 -172
rect 203 -173 204 -172
rect 204 -173 205 -172
rect 205 -173 206 -172
rect 206 -173 207 -172
rect 207 -173 208 -172
rect 208 -173 209 -172
rect 209 -173 210 -172
rect 210 -173 211 -172
rect 211 -173 212 -172
rect 212 -173 213 -172
rect 213 -173 214 -172
rect 214 -173 215 -172
rect 215 -173 216 -172
rect 216 -173 217 -172
rect 217 -173 218 -172
rect 218 -173 219 -172
rect 219 -173 220 -172
rect 220 -173 221 -172
rect 221 -173 222 -172
rect 222 -173 223 -172
rect 223 -173 224 -172
rect 224 -173 225 -172
rect 225 -173 226 -172
rect 226 -173 227 -172
rect 227 -173 228 -172
rect 228 -173 229 -172
rect 229 -173 230 -172
rect 230 -173 231 -172
rect 231 -173 232 -172
rect 232 -173 233 -172
rect 233 -173 234 -172
rect 234 -173 235 -172
rect 235 -173 236 -172
rect 236 -173 237 -172
rect 237 -173 238 -172
rect 238 -173 239 -172
rect 239 -173 240 -172
rect 240 -173 241 -172
rect 241 -173 242 -172
rect 242 -173 243 -172
rect 243 -173 244 -172
rect 244 -173 245 -172
rect 245 -173 246 -172
rect 246 -173 247 -172
rect 247 -173 248 -172
rect 248 -173 249 -172
rect 249 -173 250 -172
rect 250 -173 251 -172
rect 251 -173 252 -172
rect 252 -173 253 -172
rect 253 -173 254 -172
rect 254 -173 255 -172
rect 255 -173 256 -172
rect 256 -173 257 -172
rect 257 -173 258 -172
rect 258 -173 259 -172
rect 259 -173 260 -172
rect 260 -173 261 -172
rect 261 -173 262 -172
rect 262 -173 263 -172
rect 263 -173 264 -172
rect 264 -173 265 -172
rect 265 -173 266 -172
rect 266 -173 267 -172
rect 267 -173 268 -172
rect 268 -173 269 -172
rect 269 -173 270 -172
rect 270 -173 271 -172
rect 271 -173 272 -172
rect 272 -173 273 -172
rect 273 -173 274 -172
rect 274 -173 275 -172
rect 275 -173 276 -172
rect 276 -173 277 -172
rect 277 -173 278 -172
rect 278 -173 279 -172
rect 279 -173 280 -172
rect 280 -173 281 -172
rect 281 -173 282 -172
rect 282 -173 283 -172
rect 283 -173 284 -172
rect 284 -173 285 -172
rect 285 -173 286 -172
rect 286 -173 287 -172
rect 287 -173 288 -172
rect 288 -173 289 -172
rect 289 -173 290 -172
rect 290 -173 291 -172
rect 291 -173 292 -172
rect 292 -173 293 -172
rect 293 -173 294 -172
rect 294 -173 295 -172
rect 295 -173 296 -172
rect 296 -173 297 -172
rect 297 -173 298 -172
rect 298 -173 299 -172
rect 299 -173 300 -172
rect 300 -173 301 -172
rect 301 -173 302 -172
rect 302 -173 303 -172
rect 303 -173 304 -172
rect 304 -173 305 -172
rect 305 -173 306 -172
rect 306 -173 307 -172
rect 307 -173 308 -172
rect 308 -173 309 -172
rect 309 -173 310 -172
rect 310 -173 311 -172
rect 311 -173 312 -172
rect 312 -173 313 -172
rect 313 -173 314 -172
rect 314 -173 315 -172
rect 315 -173 316 -172
rect 316 -173 317 -172
rect 317 -173 318 -172
rect 318 -173 319 -172
rect 319 -173 320 -172
rect 320 -173 321 -172
rect 321 -173 322 -172
rect 322 -173 323 -172
rect 323 -173 324 -172
rect 324 -173 325 -172
rect 325 -173 326 -172
rect 326 -173 327 -172
rect 327 -173 328 -172
rect 328 -173 329 -172
rect 329 -173 330 -172
rect 330 -173 331 -172
rect 331 -173 332 -172
rect 332 -173 333 -172
rect 333 -173 334 -172
rect 334 -173 335 -172
rect 335 -173 336 -172
rect 336 -173 337 -172
rect 337 -173 338 -172
rect 338 -173 339 -172
rect 339 -173 340 -172
rect 340 -173 341 -172
rect 341 -173 342 -172
rect 342 -173 343 -172
rect 343 -173 344 -172
rect 344 -173 345 -172
rect 345 -173 346 -172
rect 346 -173 347 -172
rect 347 -173 348 -172
rect 348 -173 349 -172
rect 349 -173 350 -172
rect 350 -173 351 -172
rect 351 -173 352 -172
rect 352 -173 353 -172
rect 353 -173 354 -172
rect 354 -173 355 -172
rect 355 -173 356 -172
rect 356 -173 357 -172
rect 357 -173 358 -172
rect 358 -173 359 -172
rect 359 -173 360 -172
rect 360 -173 361 -172
rect 361 -173 362 -172
rect 362 -173 363 -172
rect 363 -173 364 -172
rect 364 -173 365 -172
rect 365 -173 366 -172
rect 366 -173 367 -172
rect 367 -173 368 -172
rect 368 -173 369 -172
rect 369 -173 370 -172
rect 370 -173 371 -172
rect 371 -173 372 -172
rect 372 -173 373 -172
rect 373 -173 374 -172
rect 374 -173 375 -172
rect 375 -173 376 -172
rect 376 -173 377 -172
rect 377 -173 378 -172
rect 378 -173 379 -172
rect 379 -173 380 -172
rect 380 -173 381 -172
rect 381 -173 382 -172
rect 382 -173 383 -172
rect 383 -173 384 -172
rect 384 -173 385 -172
rect 385 -173 386 -172
rect 386 -173 387 -172
rect 387 -173 388 -172
rect 388 -173 389 -172
rect 389 -173 390 -172
rect 390 -173 391 -172
rect 391 -173 392 -172
rect 392 -173 393 -172
rect 393 -173 394 -172
rect 394 -173 395 -172
rect 395 -173 396 -172
rect 396 -173 397 -172
rect 397 -173 398 -172
rect 398 -173 399 -172
rect 399 -173 400 -172
rect 400 -173 401 -172
rect 401 -173 402 -172
rect 402 -173 403 -172
rect 403 -173 404 -172
rect 404 -173 405 -172
rect 405 -173 406 -172
rect 406 -173 407 -172
rect 407 -173 408 -172
rect 408 -173 409 -172
rect 409 -173 410 -172
rect 410 -173 411 -172
rect 411 -173 412 -172
rect 412 -173 413 -172
rect 413 -173 414 -172
rect 414 -173 415 -172
rect 415 -173 416 -172
rect 416 -173 417 -172
rect 417 -173 418 -172
rect 418 -173 419 -172
rect 419 -173 420 -172
rect 420 -173 421 -172
rect 421 -173 422 -172
rect 422 -173 423 -172
rect 423 -173 424 -172
rect 424 -173 425 -172
rect 425 -173 426 -172
rect 426 -173 427 -172
rect 427 -173 428 -172
rect 428 -173 429 -172
rect 429 -173 430 -172
rect 430 -173 431 -172
rect 431 -173 432 -172
rect 432 -173 433 -172
rect 433 -173 434 -172
rect 434 -173 435 -172
rect 435 -173 436 -172
rect 436 -173 437 -172
rect 437 -173 438 -172
rect 438 -173 439 -172
rect 439 -173 440 -172
rect 440 -173 441 -172
rect 441 -173 442 -172
rect 442 -173 443 -172
rect 443 -173 444 -172
rect 444 -173 445 -172
rect 445 -173 446 -172
rect 446 -173 447 -172
rect 447 -173 448 -172
rect 448 -173 449 -172
rect 449 -173 450 -172
rect 450 -173 451 -172
rect 451 -173 452 -172
rect 452 -173 453 -172
rect 453 -173 454 -172
rect 454 -173 455 -172
rect 455 -173 456 -172
rect 456 -173 457 -172
rect 457 -173 458 -172
rect 458 -173 459 -172
rect 459 -173 460 -172
rect 460 -173 461 -172
rect 461 -173 462 -172
rect 462 -173 463 -172
rect 463 -173 464 -172
rect 464 -173 465 -172
rect 465 -173 466 -172
rect 466 -173 467 -172
rect 467 -173 468 -172
rect 468 -173 469 -172
rect 469 -173 470 -172
rect 470 -173 471 -172
rect 471 -173 472 -172
rect 472 -173 473 -172
rect 473 -173 474 -172
rect 474 -173 475 -172
rect 475 -173 476 -172
rect 476 -173 477 -172
rect 477 -173 478 -172
rect 478 -173 479 -172
rect 479 -173 480 -172
rect 2 -196 3 -195
rect 3 -196 4 -195
rect 4 -196 5 -195
rect 5 -196 6 -195
rect 6 -196 7 -195
rect 7 -196 8 -195
rect 8 -196 9 -195
rect 9 -196 10 -195
rect 10 -196 11 -195
rect 11 -196 12 -195
rect 12 -196 13 -195
rect 13 -196 14 -195
rect 14 -196 15 -195
rect 15 -196 16 -195
rect 16 -196 17 -195
rect 17 -196 18 -195
rect 18 -196 19 -195
rect 19 -196 20 -195
rect 20 -196 21 -195
rect 21 -196 22 -195
rect 22 -196 23 -195
rect 23 -196 24 -195
rect 24 -196 25 -195
rect 25 -196 26 -195
rect 26 -196 27 -195
rect 27 -196 28 -195
rect 28 -196 29 -195
rect 29 -196 30 -195
rect 30 -196 31 -195
rect 31 -196 32 -195
rect 32 -196 33 -195
rect 33 -196 34 -195
rect 34 -196 35 -195
rect 35 -196 36 -195
rect 36 -196 37 -195
rect 37 -196 38 -195
rect 38 -196 39 -195
rect 39 -196 40 -195
rect 40 -196 41 -195
rect 41 -196 42 -195
rect 42 -196 43 -195
rect 43 -196 44 -195
rect 44 -196 45 -195
rect 45 -196 46 -195
rect 46 -196 47 -195
rect 47 -196 48 -195
rect 48 -196 49 -195
rect 49 -196 50 -195
rect 50 -196 51 -195
rect 51 -196 52 -195
rect 52 -196 53 -195
rect 53 -196 54 -195
rect 54 -196 55 -195
rect 55 -196 56 -195
rect 56 -196 57 -195
rect 57 -196 58 -195
rect 58 -196 59 -195
rect 59 -196 60 -195
rect 60 -196 61 -195
rect 61 -196 62 -195
rect 62 -196 63 -195
rect 63 -196 64 -195
rect 64 -196 65 -195
rect 65 -196 66 -195
rect 66 -196 67 -195
rect 67 -196 68 -195
rect 68 -196 69 -195
rect 69 -196 70 -195
rect 70 -196 71 -195
rect 71 -196 72 -195
rect 72 -196 73 -195
rect 73 -196 74 -195
rect 74 -196 75 -195
rect 75 -196 76 -195
rect 76 -196 77 -195
rect 77 -196 78 -195
rect 78 -196 79 -195
rect 79 -196 80 -195
rect 80 -196 81 -195
rect 81 -196 82 -195
rect 82 -196 83 -195
rect 83 -196 84 -195
rect 84 -196 85 -195
rect 85 -196 86 -195
rect 86 -196 87 -195
rect 87 -196 88 -195
rect 88 -196 89 -195
rect 89 -196 90 -195
rect 90 -196 91 -195
rect 91 -196 92 -195
rect 92 -196 93 -195
rect 93 -196 94 -195
rect 94 -196 95 -195
rect 95 -196 96 -195
rect 96 -196 97 -195
rect 97 -196 98 -195
rect 98 -196 99 -195
rect 99 -196 100 -195
rect 100 -196 101 -195
rect 101 -196 102 -195
rect 102 -196 103 -195
rect 103 -196 104 -195
rect 104 -196 105 -195
rect 105 -196 106 -195
rect 106 -196 107 -195
rect 107 -196 108 -195
rect 108 -196 109 -195
rect 109 -196 110 -195
rect 110 -196 111 -195
rect 111 -196 112 -195
rect 112 -196 113 -195
rect 113 -196 114 -195
rect 114 -196 115 -195
rect 115 -196 116 -195
rect 116 -196 117 -195
rect 117 -196 118 -195
rect 118 -196 119 -195
rect 119 -196 120 -195
rect 120 -196 121 -195
rect 121 -196 122 -195
rect 122 -196 123 -195
rect 123 -196 124 -195
rect 124 -196 125 -195
rect 125 -196 126 -195
rect 126 -196 127 -195
rect 127 -196 128 -195
rect 128 -196 129 -195
rect 129 -196 130 -195
rect 130 -196 131 -195
rect 131 -196 132 -195
rect 132 -196 133 -195
rect 133 -196 134 -195
rect 134 -196 135 -195
rect 135 -196 136 -195
rect 136 -196 137 -195
rect 137 -196 138 -195
rect 138 -196 139 -195
rect 139 -196 140 -195
rect 140 -196 141 -195
rect 141 -196 142 -195
rect 142 -196 143 -195
rect 143 -196 144 -195
rect 144 -196 145 -195
rect 145 -196 146 -195
rect 146 -196 147 -195
rect 147 -196 148 -195
rect 148 -196 149 -195
rect 149 -196 150 -195
rect 150 -196 151 -195
rect 151 -196 152 -195
rect 152 -196 153 -195
rect 153 -196 154 -195
rect 154 -196 155 -195
rect 155 -196 156 -195
rect 156 -196 157 -195
rect 157 -196 158 -195
rect 158 -196 159 -195
rect 159 -196 160 -195
rect 160 -196 161 -195
rect 161 -196 162 -195
rect 162 -196 163 -195
rect 163 -196 164 -195
rect 164 -196 165 -195
rect 165 -196 166 -195
rect 166 -196 167 -195
rect 167 -196 168 -195
rect 168 -196 169 -195
rect 169 -196 170 -195
rect 170 -196 171 -195
rect 171 -196 172 -195
rect 172 -196 173 -195
rect 173 -196 174 -195
rect 174 -196 175 -195
rect 175 -196 176 -195
rect 176 -196 177 -195
rect 177 -196 178 -195
rect 178 -196 179 -195
rect 179 -196 180 -195
rect 180 -196 181 -195
rect 181 -196 182 -195
rect 182 -196 183 -195
rect 183 -196 184 -195
rect 184 -196 185 -195
rect 185 -196 186 -195
rect 186 -196 187 -195
rect 187 -196 188 -195
rect 188 -196 189 -195
rect 189 -196 190 -195
rect 190 -196 191 -195
rect 191 -196 192 -195
rect 192 -196 193 -195
rect 193 -196 194 -195
rect 194 -196 195 -195
rect 195 -196 196 -195
rect 196 -196 197 -195
rect 197 -196 198 -195
rect 198 -196 199 -195
rect 199 -196 200 -195
rect 200 -196 201 -195
rect 201 -196 202 -195
rect 202 -196 203 -195
rect 203 -196 204 -195
rect 204 -196 205 -195
rect 205 -196 206 -195
rect 206 -196 207 -195
rect 207 -196 208 -195
rect 208 -196 209 -195
rect 209 -196 210 -195
rect 210 -196 211 -195
rect 211 -196 212 -195
rect 212 -196 213 -195
rect 213 -196 214 -195
rect 214 -196 215 -195
rect 215 -196 216 -195
rect 216 -196 217 -195
rect 217 -196 218 -195
rect 218 -196 219 -195
rect 219 -196 220 -195
rect 220 -196 221 -195
rect 221 -196 222 -195
rect 222 -196 223 -195
rect 223 -196 224 -195
rect 224 -196 225 -195
rect 225 -196 226 -195
rect 226 -196 227 -195
rect 227 -196 228 -195
rect 228 -196 229 -195
rect 229 -196 230 -195
rect 230 -196 231 -195
rect 231 -196 232 -195
rect 232 -196 233 -195
rect 233 -196 234 -195
rect 234 -196 235 -195
rect 235 -196 236 -195
rect 236 -196 237 -195
rect 237 -196 238 -195
rect 238 -196 239 -195
rect 239 -196 240 -195
rect 240 -196 241 -195
rect 241 -196 242 -195
rect 242 -196 243 -195
rect 243 -196 244 -195
rect 244 -196 245 -195
rect 245 -196 246 -195
rect 246 -196 247 -195
rect 247 -196 248 -195
rect 248 -196 249 -195
rect 249 -196 250 -195
rect 250 -196 251 -195
rect 251 -196 252 -195
rect 252 -196 253 -195
rect 253 -196 254 -195
rect 254 -196 255 -195
rect 255 -196 256 -195
rect 256 -196 257 -195
rect 257 -196 258 -195
rect 258 -196 259 -195
rect 259 -196 260 -195
rect 260 -196 261 -195
rect 261 -196 262 -195
rect 262 -196 263 -195
rect 263 -196 264 -195
rect 264 -196 265 -195
rect 265 -196 266 -195
rect 266 -196 267 -195
rect 267 -196 268 -195
rect 268 -196 269 -195
rect 269 -196 270 -195
rect 270 -196 271 -195
rect 271 -196 272 -195
rect 272 -196 273 -195
rect 273 -196 274 -195
rect 274 -196 275 -195
rect 275 -196 276 -195
rect 276 -196 277 -195
rect 277 -196 278 -195
rect 278 -196 279 -195
rect 279 -196 280 -195
rect 280 -196 281 -195
rect 281 -196 282 -195
rect 282 -196 283 -195
rect 283 -196 284 -195
rect 284 -196 285 -195
rect 285 -196 286 -195
rect 286 -196 287 -195
rect 287 -196 288 -195
rect 288 -196 289 -195
rect 289 -196 290 -195
rect 290 -196 291 -195
rect 291 -196 292 -195
rect 292 -196 293 -195
rect 293 -196 294 -195
rect 294 -196 295 -195
rect 295 -196 296 -195
rect 296 -196 297 -195
rect 297 -196 298 -195
rect 298 -196 299 -195
rect 299 -196 300 -195
rect 300 -196 301 -195
rect 301 -196 302 -195
rect 302 -196 303 -195
rect 303 -196 304 -195
rect 304 -196 305 -195
rect 305 -196 306 -195
rect 306 -196 307 -195
rect 307 -196 308 -195
rect 308 -196 309 -195
rect 309 -196 310 -195
rect 310 -196 311 -195
rect 311 -196 312 -195
rect 312 -196 313 -195
rect 313 -196 314 -195
rect 314 -196 315 -195
rect 315 -196 316 -195
rect 316 -196 317 -195
rect 317 -196 318 -195
rect 318 -196 319 -195
rect 319 -196 320 -195
rect 320 -196 321 -195
rect 321 -196 322 -195
rect 322 -196 323 -195
rect 323 -196 324 -195
rect 324 -196 325 -195
rect 325 -196 326 -195
rect 326 -196 327 -195
rect 327 -196 328 -195
rect 328 -196 329 -195
rect 329 -196 330 -195
rect 330 -196 331 -195
rect 331 -196 332 -195
rect 332 -196 333 -195
rect 333 -196 334 -195
rect 334 -196 335 -195
rect 335 -196 336 -195
rect 336 -196 337 -195
rect 337 -196 338 -195
rect 338 -196 339 -195
rect 339 -196 340 -195
rect 340 -196 341 -195
rect 341 -196 342 -195
rect 342 -196 343 -195
rect 343 -196 344 -195
rect 344 -196 345 -195
rect 345 -196 346 -195
rect 346 -196 347 -195
rect 347 -196 348 -195
rect 348 -196 349 -195
rect 349 -196 350 -195
rect 350 -196 351 -195
rect 351 -196 352 -195
rect 352 -196 353 -195
rect 353 -196 354 -195
rect 354 -196 355 -195
rect 355 -196 356 -195
rect 356 -196 357 -195
rect 357 -196 358 -195
rect 358 -196 359 -195
rect 359 -196 360 -195
rect 360 -196 361 -195
rect 361 -196 362 -195
rect 362 -196 363 -195
rect 363 -196 364 -195
rect 364 -196 365 -195
rect 365 -196 366 -195
rect 366 -196 367 -195
rect 367 -196 368 -195
rect 368 -196 369 -195
rect 369 -196 370 -195
rect 370 -196 371 -195
rect 371 -196 372 -195
rect 372 -196 373 -195
rect 373 -196 374 -195
rect 374 -196 375 -195
rect 375 -196 376 -195
rect 376 -196 377 -195
rect 377 -196 378 -195
rect 378 -196 379 -195
rect 379 -196 380 -195
rect 380 -196 381 -195
rect 381 -196 382 -195
rect 382 -196 383 -195
rect 383 -196 384 -195
rect 384 -196 385 -195
rect 385 -196 386 -195
rect 386 -196 387 -195
rect 387 -196 388 -195
rect 388 -196 389 -195
rect 389 -196 390 -195
rect 390 -196 391 -195
rect 391 -196 392 -195
rect 392 -196 393 -195
rect 393 -196 394 -195
rect 394 -196 395 -195
rect 395 -196 396 -195
rect 396 -196 397 -195
rect 397 -196 398 -195
rect 398 -196 399 -195
rect 399 -196 400 -195
rect 400 -196 401 -195
rect 401 -196 402 -195
rect 402 -196 403 -195
rect 403 -196 404 -195
rect 404 -196 405 -195
rect 405 -196 406 -195
rect 406 -196 407 -195
rect 407 -196 408 -195
rect 408 -196 409 -195
rect 409 -196 410 -195
rect 410 -196 411 -195
rect 411 -196 412 -195
rect 412 -196 413 -195
rect 413 -196 414 -195
rect 414 -196 415 -195
rect 415 -196 416 -195
rect 416 -196 417 -195
rect 417 -196 418 -195
rect 418 -196 419 -195
rect 419 -196 420 -195
rect 420 -196 421 -195
rect 421 -196 422 -195
rect 422 -196 423 -195
rect 423 -196 424 -195
rect 424 -196 425 -195
rect 425 -196 426 -195
rect 426 -196 427 -195
rect 427 -196 428 -195
rect 428 -196 429 -195
rect 429 -196 430 -195
rect 430 -196 431 -195
rect 431 -196 432 -195
rect 432 -196 433 -195
rect 433 -196 434 -195
rect 434 -196 435 -195
rect 435 -196 436 -195
rect 436 -196 437 -195
rect 437 -196 438 -195
rect 438 -196 439 -195
rect 439 -196 440 -195
rect 440 -196 441 -195
rect 441 -196 442 -195
rect 442 -196 443 -195
rect 443 -196 444 -195
rect 444 -196 445 -195
rect 445 -196 446 -195
rect 446 -196 447 -195
rect 447 -196 448 -195
rect 448 -196 449 -195
rect 449 -196 450 -195
rect 450 -196 451 -195
rect 451 -196 452 -195
rect 452 -196 453 -195
rect 453 -196 454 -195
rect 454 -196 455 -195
rect 455 -196 456 -195
rect 456 -196 457 -195
rect 457 -196 458 -195
rect 458 -196 459 -195
rect 459 -196 460 -195
rect 460 -196 461 -195
rect 461 -196 462 -195
rect 462 -196 463 -195
rect 463 -196 464 -195
rect 464 -196 465 -195
rect 465 -196 466 -195
rect 466 -196 467 -195
rect 467 -196 468 -195
rect 468 -196 469 -195
rect 469 -196 470 -195
rect 470 -196 471 -195
rect 471 -196 472 -195
rect 472 -196 473 -195
rect 473 -196 474 -195
rect 474 -196 475 -195
rect 475 -196 476 -195
rect 476 -196 477 -195
rect 477 -196 478 -195
rect 478 -196 479 -195
rect 479 -196 480 -195
rect 2 -197 3 -196
rect 3 -197 4 -196
rect 4 -197 5 -196
rect 5 -197 6 -196
rect 6 -197 7 -196
rect 7 -197 8 -196
rect 8 -197 9 -196
rect 9 -197 10 -196
rect 10 -197 11 -196
rect 11 -197 12 -196
rect 12 -197 13 -196
rect 13 -197 14 -196
rect 14 -197 15 -196
rect 15 -197 16 -196
rect 16 -197 17 -196
rect 17 -197 18 -196
rect 18 -197 19 -196
rect 19 -197 20 -196
rect 20 -197 21 -196
rect 21 -197 22 -196
rect 22 -197 23 -196
rect 23 -197 24 -196
rect 24 -197 25 -196
rect 25 -197 26 -196
rect 26 -197 27 -196
rect 27 -197 28 -196
rect 28 -197 29 -196
rect 29 -197 30 -196
rect 30 -197 31 -196
rect 31 -197 32 -196
rect 32 -197 33 -196
rect 33 -197 34 -196
rect 34 -197 35 -196
rect 35 -197 36 -196
rect 36 -197 37 -196
rect 37 -197 38 -196
rect 38 -197 39 -196
rect 39 -197 40 -196
rect 40 -197 41 -196
rect 41 -197 42 -196
rect 42 -197 43 -196
rect 43 -197 44 -196
rect 44 -197 45 -196
rect 45 -197 46 -196
rect 46 -197 47 -196
rect 47 -197 48 -196
rect 48 -197 49 -196
rect 49 -197 50 -196
rect 50 -197 51 -196
rect 51 -197 52 -196
rect 52 -197 53 -196
rect 53 -197 54 -196
rect 54 -197 55 -196
rect 55 -197 56 -196
rect 56 -197 57 -196
rect 57 -197 58 -196
rect 58 -197 59 -196
rect 59 -197 60 -196
rect 60 -197 61 -196
rect 61 -197 62 -196
rect 62 -197 63 -196
rect 63 -197 64 -196
rect 64 -197 65 -196
rect 65 -197 66 -196
rect 66 -197 67 -196
rect 67 -197 68 -196
rect 68 -197 69 -196
rect 69 -197 70 -196
rect 70 -197 71 -196
rect 71 -197 72 -196
rect 72 -197 73 -196
rect 73 -197 74 -196
rect 74 -197 75 -196
rect 75 -197 76 -196
rect 76 -197 77 -196
rect 77 -197 78 -196
rect 78 -197 79 -196
rect 79 -197 80 -196
rect 80 -197 81 -196
rect 81 -197 82 -196
rect 82 -197 83 -196
rect 83 -197 84 -196
rect 84 -197 85 -196
rect 85 -197 86 -196
rect 86 -197 87 -196
rect 87 -197 88 -196
rect 88 -197 89 -196
rect 89 -197 90 -196
rect 90 -197 91 -196
rect 91 -197 92 -196
rect 92 -197 93 -196
rect 93 -197 94 -196
rect 94 -197 95 -196
rect 95 -197 96 -196
rect 96 -197 97 -196
rect 97 -197 98 -196
rect 98 -197 99 -196
rect 99 -197 100 -196
rect 100 -197 101 -196
rect 101 -197 102 -196
rect 102 -197 103 -196
rect 103 -197 104 -196
rect 104 -197 105 -196
rect 105 -197 106 -196
rect 106 -197 107 -196
rect 107 -197 108 -196
rect 108 -197 109 -196
rect 109 -197 110 -196
rect 110 -197 111 -196
rect 111 -197 112 -196
rect 112 -197 113 -196
rect 113 -197 114 -196
rect 114 -197 115 -196
rect 115 -197 116 -196
rect 116 -197 117 -196
rect 117 -197 118 -196
rect 118 -197 119 -196
rect 119 -197 120 -196
rect 120 -197 121 -196
rect 121 -197 122 -196
rect 122 -197 123 -196
rect 123 -197 124 -196
rect 124 -197 125 -196
rect 125 -197 126 -196
rect 126 -197 127 -196
rect 127 -197 128 -196
rect 128 -197 129 -196
rect 129 -197 130 -196
rect 130 -197 131 -196
rect 131 -197 132 -196
rect 132 -197 133 -196
rect 133 -197 134 -196
rect 134 -197 135 -196
rect 135 -197 136 -196
rect 136 -197 137 -196
rect 137 -197 138 -196
rect 138 -197 139 -196
rect 139 -197 140 -196
rect 140 -197 141 -196
rect 141 -197 142 -196
rect 142 -197 143 -196
rect 143 -197 144 -196
rect 144 -197 145 -196
rect 145 -197 146 -196
rect 146 -197 147 -196
rect 147 -197 148 -196
rect 148 -197 149 -196
rect 149 -197 150 -196
rect 150 -197 151 -196
rect 151 -197 152 -196
rect 152 -197 153 -196
rect 153 -197 154 -196
rect 154 -197 155 -196
rect 155 -197 156 -196
rect 156 -197 157 -196
rect 157 -197 158 -196
rect 158 -197 159 -196
rect 159 -197 160 -196
rect 160 -197 161 -196
rect 161 -197 162 -196
rect 162 -197 163 -196
rect 163 -197 164 -196
rect 164 -197 165 -196
rect 165 -197 166 -196
rect 166 -197 167 -196
rect 167 -197 168 -196
rect 168 -197 169 -196
rect 169 -197 170 -196
rect 170 -197 171 -196
rect 171 -197 172 -196
rect 172 -197 173 -196
rect 173 -197 174 -196
rect 174 -197 175 -196
rect 175 -197 176 -196
rect 176 -197 177 -196
rect 177 -197 178 -196
rect 178 -197 179 -196
rect 179 -197 180 -196
rect 180 -197 181 -196
rect 181 -197 182 -196
rect 182 -197 183 -196
rect 183 -197 184 -196
rect 184 -197 185 -196
rect 185 -197 186 -196
rect 186 -197 187 -196
rect 187 -197 188 -196
rect 188 -197 189 -196
rect 189 -197 190 -196
rect 190 -197 191 -196
rect 191 -197 192 -196
rect 192 -197 193 -196
rect 193 -197 194 -196
rect 194 -197 195 -196
rect 195 -197 196 -196
rect 196 -197 197 -196
rect 197 -197 198 -196
rect 198 -197 199 -196
rect 199 -197 200 -196
rect 200 -197 201 -196
rect 201 -197 202 -196
rect 202 -197 203 -196
rect 203 -197 204 -196
rect 204 -197 205 -196
rect 205 -197 206 -196
rect 206 -197 207 -196
rect 207 -197 208 -196
rect 208 -197 209 -196
rect 209 -197 210 -196
rect 210 -197 211 -196
rect 211 -197 212 -196
rect 212 -197 213 -196
rect 213 -197 214 -196
rect 214 -197 215 -196
rect 215 -197 216 -196
rect 216 -197 217 -196
rect 217 -197 218 -196
rect 218 -197 219 -196
rect 219 -197 220 -196
rect 220 -197 221 -196
rect 221 -197 222 -196
rect 222 -197 223 -196
rect 223 -197 224 -196
rect 224 -197 225 -196
rect 225 -197 226 -196
rect 226 -197 227 -196
rect 227 -197 228 -196
rect 228 -197 229 -196
rect 229 -197 230 -196
rect 230 -197 231 -196
rect 231 -197 232 -196
rect 232 -197 233 -196
rect 233 -197 234 -196
rect 234 -197 235 -196
rect 235 -197 236 -196
rect 236 -197 237 -196
rect 237 -197 238 -196
rect 238 -197 239 -196
rect 239 -197 240 -196
rect 240 -197 241 -196
rect 241 -197 242 -196
rect 242 -197 243 -196
rect 243 -197 244 -196
rect 244 -197 245 -196
rect 245 -197 246 -196
rect 246 -197 247 -196
rect 247 -197 248 -196
rect 248 -197 249 -196
rect 249 -197 250 -196
rect 250 -197 251 -196
rect 251 -197 252 -196
rect 252 -197 253 -196
rect 253 -197 254 -196
rect 254 -197 255 -196
rect 255 -197 256 -196
rect 256 -197 257 -196
rect 257 -197 258 -196
rect 258 -197 259 -196
rect 259 -197 260 -196
rect 260 -197 261 -196
rect 261 -197 262 -196
rect 262 -197 263 -196
rect 263 -197 264 -196
rect 264 -197 265 -196
rect 265 -197 266 -196
rect 266 -197 267 -196
rect 267 -197 268 -196
rect 268 -197 269 -196
rect 269 -197 270 -196
rect 270 -197 271 -196
rect 271 -197 272 -196
rect 272 -197 273 -196
rect 273 -197 274 -196
rect 274 -197 275 -196
rect 275 -197 276 -196
rect 276 -197 277 -196
rect 277 -197 278 -196
rect 278 -197 279 -196
rect 279 -197 280 -196
rect 280 -197 281 -196
rect 281 -197 282 -196
rect 282 -197 283 -196
rect 283 -197 284 -196
rect 284 -197 285 -196
rect 285 -197 286 -196
rect 286 -197 287 -196
rect 287 -197 288 -196
rect 288 -197 289 -196
rect 289 -197 290 -196
rect 290 -197 291 -196
rect 291 -197 292 -196
rect 292 -197 293 -196
rect 293 -197 294 -196
rect 294 -197 295 -196
rect 295 -197 296 -196
rect 296 -197 297 -196
rect 297 -197 298 -196
rect 298 -197 299 -196
rect 299 -197 300 -196
rect 300 -197 301 -196
rect 301 -197 302 -196
rect 302 -197 303 -196
rect 303 -197 304 -196
rect 304 -197 305 -196
rect 305 -197 306 -196
rect 306 -197 307 -196
rect 307 -197 308 -196
rect 308 -197 309 -196
rect 309 -197 310 -196
rect 310 -197 311 -196
rect 311 -197 312 -196
rect 312 -197 313 -196
rect 313 -197 314 -196
rect 314 -197 315 -196
rect 315 -197 316 -196
rect 316 -197 317 -196
rect 317 -197 318 -196
rect 318 -197 319 -196
rect 319 -197 320 -196
rect 320 -197 321 -196
rect 321 -197 322 -196
rect 322 -197 323 -196
rect 323 -197 324 -196
rect 324 -197 325 -196
rect 325 -197 326 -196
rect 326 -197 327 -196
rect 327 -197 328 -196
rect 328 -197 329 -196
rect 329 -197 330 -196
rect 330 -197 331 -196
rect 331 -197 332 -196
rect 332 -197 333 -196
rect 333 -197 334 -196
rect 334 -197 335 -196
rect 335 -197 336 -196
rect 336 -197 337 -196
rect 337 -197 338 -196
rect 338 -197 339 -196
rect 339 -197 340 -196
rect 340 -197 341 -196
rect 341 -197 342 -196
rect 342 -197 343 -196
rect 343 -197 344 -196
rect 344 -197 345 -196
rect 345 -197 346 -196
rect 346 -197 347 -196
rect 347 -197 348 -196
rect 348 -197 349 -196
rect 349 -197 350 -196
rect 350 -197 351 -196
rect 351 -197 352 -196
rect 352 -197 353 -196
rect 353 -197 354 -196
rect 354 -197 355 -196
rect 355 -197 356 -196
rect 356 -197 357 -196
rect 357 -197 358 -196
rect 358 -197 359 -196
rect 359 -197 360 -196
rect 360 -197 361 -196
rect 361 -197 362 -196
rect 362 -197 363 -196
rect 363 -197 364 -196
rect 364 -197 365 -196
rect 365 -197 366 -196
rect 366 -197 367 -196
rect 367 -197 368 -196
rect 368 -197 369 -196
rect 369 -197 370 -196
rect 370 -197 371 -196
rect 371 -197 372 -196
rect 372 -197 373 -196
rect 373 -197 374 -196
rect 374 -197 375 -196
rect 375 -197 376 -196
rect 376 -197 377 -196
rect 377 -197 378 -196
rect 378 -197 379 -196
rect 379 -197 380 -196
rect 380 -197 381 -196
rect 381 -197 382 -196
rect 382 -197 383 -196
rect 383 -197 384 -196
rect 384 -197 385 -196
rect 385 -197 386 -196
rect 386 -197 387 -196
rect 387 -197 388 -196
rect 388 -197 389 -196
rect 389 -197 390 -196
rect 390 -197 391 -196
rect 391 -197 392 -196
rect 392 -197 393 -196
rect 393 -197 394 -196
rect 394 -197 395 -196
rect 395 -197 396 -196
rect 396 -197 397 -196
rect 397 -197 398 -196
rect 398 -197 399 -196
rect 399 -197 400 -196
rect 400 -197 401 -196
rect 401 -197 402 -196
rect 402 -197 403 -196
rect 403 -197 404 -196
rect 404 -197 405 -196
rect 405 -197 406 -196
rect 406 -197 407 -196
rect 407 -197 408 -196
rect 408 -197 409 -196
rect 409 -197 410 -196
rect 410 -197 411 -196
rect 411 -197 412 -196
rect 412 -197 413 -196
rect 413 -197 414 -196
rect 414 -197 415 -196
rect 415 -197 416 -196
rect 416 -197 417 -196
rect 417 -197 418 -196
rect 418 -197 419 -196
rect 419 -197 420 -196
rect 420 -197 421 -196
rect 421 -197 422 -196
rect 422 -197 423 -196
rect 423 -197 424 -196
rect 424 -197 425 -196
rect 425 -197 426 -196
rect 426 -197 427 -196
rect 427 -197 428 -196
rect 428 -197 429 -196
rect 429 -197 430 -196
rect 430 -197 431 -196
rect 431 -197 432 -196
rect 432 -197 433 -196
rect 433 -197 434 -196
rect 434 -197 435 -196
rect 435 -197 436 -196
rect 436 -197 437 -196
rect 437 -197 438 -196
rect 438 -197 439 -196
rect 439 -197 440 -196
rect 440 -197 441 -196
rect 441 -197 442 -196
rect 442 -197 443 -196
rect 443 -197 444 -196
rect 444 -197 445 -196
rect 445 -197 446 -196
rect 446 -197 447 -196
rect 447 -197 448 -196
rect 448 -197 449 -196
rect 449 -197 450 -196
rect 450 -197 451 -196
rect 451 -197 452 -196
rect 452 -197 453 -196
rect 453 -197 454 -196
rect 454 -197 455 -196
rect 455 -197 456 -196
rect 456 -197 457 -196
rect 457 -197 458 -196
rect 458 -197 459 -196
rect 459 -197 460 -196
rect 460 -197 461 -196
rect 461 -197 462 -196
rect 462 -197 463 -196
rect 463 -197 464 -196
rect 464 -197 465 -196
rect 465 -197 466 -196
rect 466 -197 467 -196
rect 467 -197 468 -196
rect 468 -197 469 -196
rect 469 -197 470 -196
rect 470 -197 471 -196
rect 471 -197 472 -196
rect 472 -197 473 -196
rect 473 -197 474 -196
rect 474 -197 475 -196
rect 475 -197 476 -196
rect 476 -197 477 -196
rect 477 -197 478 -196
rect 478 -197 479 -196
rect 479 -197 480 -196
rect 2 -198 3 -197
rect 3 -198 4 -197
rect 4 -198 5 -197
rect 5 -198 6 -197
rect 6 -198 7 -197
rect 7 -198 8 -197
rect 8 -198 9 -197
rect 9 -198 10 -197
rect 10 -198 11 -197
rect 11 -198 12 -197
rect 12 -198 13 -197
rect 13 -198 14 -197
rect 14 -198 15 -197
rect 15 -198 16 -197
rect 16 -198 17 -197
rect 17 -198 18 -197
rect 18 -198 19 -197
rect 19 -198 20 -197
rect 20 -198 21 -197
rect 21 -198 22 -197
rect 22 -198 23 -197
rect 23 -198 24 -197
rect 24 -198 25 -197
rect 25 -198 26 -197
rect 26 -198 27 -197
rect 27 -198 28 -197
rect 28 -198 29 -197
rect 29 -198 30 -197
rect 30 -198 31 -197
rect 31 -198 32 -197
rect 32 -198 33 -197
rect 33 -198 34 -197
rect 34 -198 35 -197
rect 35 -198 36 -197
rect 36 -198 37 -197
rect 37 -198 38 -197
rect 38 -198 39 -197
rect 39 -198 40 -197
rect 40 -198 41 -197
rect 41 -198 42 -197
rect 42 -198 43 -197
rect 43 -198 44 -197
rect 44 -198 45 -197
rect 45 -198 46 -197
rect 46 -198 47 -197
rect 47 -198 48 -197
rect 48 -198 49 -197
rect 49 -198 50 -197
rect 50 -198 51 -197
rect 51 -198 52 -197
rect 52 -198 53 -197
rect 53 -198 54 -197
rect 54 -198 55 -197
rect 55 -198 56 -197
rect 56 -198 57 -197
rect 57 -198 58 -197
rect 58 -198 59 -197
rect 59 -198 60 -197
rect 60 -198 61 -197
rect 61 -198 62 -197
rect 62 -198 63 -197
rect 63 -198 64 -197
rect 64 -198 65 -197
rect 65 -198 66 -197
rect 66 -198 67 -197
rect 67 -198 68 -197
rect 68 -198 69 -197
rect 69 -198 70 -197
rect 70 -198 71 -197
rect 71 -198 72 -197
rect 72 -198 73 -197
rect 73 -198 74 -197
rect 74 -198 75 -197
rect 75 -198 76 -197
rect 76 -198 77 -197
rect 77 -198 78 -197
rect 78 -198 79 -197
rect 79 -198 80 -197
rect 80 -198 81 -197
rect 81 -198 82 -197
rect 82 -198 83 -197
rect 83 -198 84 -197
rect 84 -198 85 -197
rect 85 -198 86 -197
rect 86 -198 87 -197
rect 87 -198 88 -197
rect 88 -198 89 -197
rect 89 -198 90 -197
rect 90 -198 91 -197
rect 91 -198 92 -197
rect 92 -198 93 -197
rect 93 -198 94 -197
rect 94 -198 95 -197
rect 95 -198 96 -197
rect 96 -198 97 -197
rect 97 -198 98 -197
rect 98 -198 99 -197
rect 99 -198 100 -197
rect 100 -198 101 -197
rect 101 -198 102 -197
rect 102 -198 103 -197
rect 103 -198 104 -197
rect 104 -198 105 -197
rect 105 -198 106 -197
rect 106 -198 107 -197
rect 107 -198 108 -197
rect 108 -198 109 -197
rect 109 -198 110 -197
rect 110 -198 111 -197
rect 111 -198 112 -197
rect 112 -198 113 -197
rect 113 -198 114 -197
rect 114 -198 115 -197
rect 115 -198 116 -197
rect 116 -198 117 -197
rect 117 -198 118 -197
rect 118 -198 119 -197
rect 119 -198 120 -197
rect 120 -198 121 -197
rect 121 -198 122 -197
rect 122 -198 123 -197
rect 123 -198 124 -197
rect 124 -198 125 -197
rect 125 -198 126 -197
rect 126 -198 127 -197
rect 127 -198 128 -197
rect 128 -198 129 -197
rect 129 -198 130 -197
rect 130 -198 131 -197
rect 131 -198 132 -197
rect 132 -198 133 -197
rect 133 -198 134 -197
rect 134 -198 135 -197
rect 135 -198 136 -197
rect 136 -198 137 -197
rect 137 -198 138 -197
rect 138 -198 139 -197
rect 139 -198 140 -197
rect 140 -198 141 -197
rect 141 -198 142 -197
rect 142 -198 143 -197
rect 143 -198 144 -197
rect 144 -198 145 -197
rect 145 -198 146 -197
rect 146 -198 147 -197
rect 147 -198 148 -197
rect 148 -198 149 -197
rect 149 -198 150 -197
rect 150 -198 151 -197
rect 151 -198 152 -197
rect 152 -198 153 -197
rect 153 -198 154 -197
rect 154 -198 155 -197
rect 155 -198 156 -197
rect 156 -198 157 -197
rect 157 -198 158 -197
rect 158 -198 159 -197
rect 159 -198 160 -197
rect 160 -198 161 -197
rect 161 -198 162 -197
rect 162 -198 163 -197
rect 163 -198 164 -197
rect 164 -198 165 -197
rect 165 -198 166 -197
rect 166 -198 167 -197
rect 167 -198 168 -197
rect 168 -198 169 -197
rect 169 -198 170 -197
rect 170 -198 171 -197
rect 171 -198 172 -197
rect 172 -198 173 -197
rect 173 -198 174 -197
rect 174 -198 175 -197
rect 175 -198 176 -197
rect 176 -198 177 -197
rect 177 -198 178 -197
rect 178 -198 179 -197
rect 179 -198 180 -197
rect 180 -198 181 -197
rect 181 -198 182 -197
rect 182 -198 183 -197
rect 183 -198 184 -197
rect 184 -198 185 -197
rect 185 -198 186 -197
rect 186 -198 187 -197
rect 187 -198 188 -197
rect 188 -198 189 -197
rect 189 -198 190 -197
rect 190 -198 191 -197
rect 191 -198 192 -197
rect 192 -198 193 -197
rect 193 -198 194 -197
rect 194 -198 195 -197
rect 195 -198 196 -197
rect 196 -198 197 -197
rect 197 -198 198 -197
rect 198 -198 199 -197
rect 199 -198 200 -197
rect 200 -198 201 -197
rect 201 -198 202 -197
rect 202 -198 203 -197
rect 203 -198 204 -197
rect 204 -198 205 -197
rect 205 -198 206 -197
rect 206 -198 207 -197
rect 207 -198 208 -197
rect 208 -198 209 -197
rect 209 -198 210 -197
rect 210 -198 211 -197
rect 211 -198 212 -197
rect 212 -198 213 -197
rect 213 -198 214 -197
rect 214 -198 215 -197
rect 215 -198 216 -197
rect 216 -198 217 -197
rect 217 -198 218 -197
rect 218 -198 219 -197
rect 219 -198 220 -197
rect 220 -198 221 -197
rect 221 -198 222 -197
rect 222 -198 223 -197
rect 223 -198 224 -197
rect 224 -198 225 -197
rect 225 -198 226 -197
rect 226 -198 227 -197
rect 227 -198 228 -197
rect 228 -198 229 -197
rect 229 -198 230 -197
rect 230 -198 231 -197
rect 231 -198 232 -197
rect 232 -198 233 -197
rect 233 -198 234 -197
rect 234 -198 235 -197
rect 235 -198 236 -197
rect 236 -198 237 -197
rect 237 -198 238 -197
rect 238 -198 239 -197
rect 239 -198 240 -197
rect 240 -198 241 -197
rect 241 -198 242 -197
rect 242 -198 243 -197
rect 243 -198 244 -197
rect 244 -198 245 -197
rect 245 -198 246 -197
rect 246 -198 247 -197
rect 247 -198 248 -197
rect 248 -198 249 -197
rect 249 -198 250 -197
rect 250 -198 251 -197
rect 251 -198 252 -197
rect 252 -198 253 -197
rect 253 -198 254 -197
rect 254 -198 255 -197
rect 255 -198 256 -197
rect 256 -198 257 -197
rect 257 -198 258 -197
rect 258 -198 259 -197
rect 259 -198 260 -197
rect 260 -198 261 -197
rect 261 -198 262 -197
rect 262 -198 263 -197
rect 263 -198 264 -197
rect 264 -198 265 -197
rect 265 -198 266 -197
rect 266 -198 267 -197
rect 267 -198 268 -197
rect 268 -198 269 -197
rect 269 -198 270 -197
rect 270 -198 271 -197
rect 271 -198 272 -197
rect 272 -198 273 -197
rect 273 -198 274 -197
rect 274 -198 275 -197
rect 275 -198 276 -197
rect 276 -198 277 -197
rect 277 -198 278 -197
rect 278 -198 279 -197
rect 279 -198 280 -197
rect 280 -198 281 -197
rect 281 -198 282 -197
rect 282 -198 283 -197
rect 283 -198 284 -197
rect 284 -198 285 -197
rect 285 -198 286 -197
rect 286 -198 287 -197
rect 287 -198 288 -197
rect 288 -198 289 -197
rect 289 -198 290 -197
rect 290 -198 291 -197
rect 291 -198 292 -197
rect 292 -198 293 -197
rect 293 -198 294 -197
rect 294 -198 295 -197
rect 295 -198 296 -197
rect 296 -198 297 -197
rect 297 -198 298 -197
rect 298 -198 299 -197
rect 299 -198 300 -197
rect 300 -198 301 -197
rect 301 -198 302 -197
rect 302 -198 303 -197
rect 303 -198 304 -197
rect 304 -198 305 -197
rect 305 -198 306 -197
rect 306 -198 307 -197
rect 307 -198 308 -197
rect 308 -198 309 -197
rect 309 -198 310 -197
rect 310 -198 311 -197
rect 311 -198 312 -197
rect 312 -198 313 -197
rect 313 -198 314 -197
rect 314 -198 315 -197
rect 315 -198 316 -197
rect 316 -198 317 -197
rect 317 -198 318 -197
rect 318 -198 319 -197
rect 319 -198 320 -197
rect 320 -198 321 -197
rect 321 -198 322 -197
rect 322 -198 323 -197
rect 323 -198 324 -197
rect 324 -198 325 -197
rect 325 -198 326 -197
rect 326 -198 327 -197
rect 327 -198 328 -197
rect 328 -198 329 -197
rect 329 -198 330 -197
rect 330 -198 331 -197
rect 331 -198 332 -197
rect 332 -198 333 -197
rect 333 -198 334 -197
rect 334 -198 335 -197
rect 335 -198 336 -197
rect 336 -198 337 -197
rect 337 -198 338 -197
rect 338 -198 339 -197
rect 339 -198 340 -197
rect 340 -198 341 -197
rect 341 -198 342 -197
rect 342 -198 343 -197
rect 343 -198 344 -197
rect 344 -198 345 -197
rect 345 -198 346 -197
rect 346 -198 347 -197
rect 347 -198 348 -197
rect 348 -198 349 -197
rect 349 -198 350 -197
rect 350 -198 351 -197
rect 351 -198 352 -197
rect 352 -198 353 -197
rect 353 -198 354 -197
rect 354 -198 355 -197
rect 355 -198 356 -197
rect 356 -198 357 -197
rect 357 -198 358 -197
rect 358 -198 359 -197
rect 359 -198 360 -197
rect 360 -198 361 -197
rect 361 -198 362 -197
rect 362 -198 363 -197
rect 363 -198 364 -197
rect 364 -198 365 -197
rect 365 -198 366 -197
rect 366 -198 367 -197
rect 367 -198 368 -197
rect 368 -198 369 -197
rect 369 -198 370 -197
rect 370 -198 371 -197
rect 371 -198 372 -197
rect 372 -198 373 -197
rect 373 -198 374 -197
rect 374 -198 375 -197
rect 375 -198 376 -197
rect 376 -198 377 -197
rect 377 -198 378 -197
rect 378 -198 379 -197
rect 379 -198 380 -197
rect 380 -198 381 -197
rect 381 -198 382 -197
rect 382 -198 383 -197
rect 383 -198 384 -197
rect 384 -198 385 -197
rect 385 -198 386 -197
rect 386 -198 387 -197
rect 387 -198 388 -197
rect 388 -198 389 -197
rect 389 -198 390 -197
rect 390 -198 391 -197
rect 391 -198 392 -197
rect 392 -198 393 -197
rect 393 -198 394 -197
rect 394 -198 395 -197
rect 395 -198 396 -197
rect 396 -198 397 -197
rect 397 -198 398 -197
rect 398 -198 399 -197
rect 399 -198 400 -197
rect 400 -198 401 -197
rect 401 -198 402 -197
rect 402 -198 403 -197
rect 403 -198 404 -197
rect 404 -198 405 -197
rect 405 -198 406 -197
rect 406 -198 407 -197
rect 407 -198 408 -197
rect 408 -198 409 -197
rect 409 -198 410 -197
rect 410 -198 411 -197
rect 411 -198 412 -197
rect 412 -198 413 -197
rect 413 -198 414 -197
rect 414 -198 415 -197
rect 415 -198 416 -197
rect 416 -198 417 -197
rect 417 -198 418 -197
rect 418 -198 419 -197
rect 419 -198 420 -197
rect 420 -198 421 -197
rect 421 -198 422 -197
rect 422 -198 423 -197
rect 423 -198 424 -197
rect 424 -198 425 -197
rect 425 -198 426 -197
rect 426 -198 427 -197
rect 427 -198 428 -197
rect 428 -198 429 -197
rect 429 -198 430 -197
rect 430 -198 431 -197
rect 431 -198 432 -197
rect 432 -198 433 -197
rect 433 -198 434 -197
rect 434 -198 435 -197
rect 435 -198 436 -197
rect 436 -198 437 -197
rect 437 -198 438 -197
rect 438 -198 439 -197
rect 439 -198 440 -197
rect 440 -198 441 -197
rect 441 -198 442 -197
rect 442 -198 443 -197
rect 443 -198 444 -197
rect 444 -198 445 -197
rect 445 -198 446 -197
rect 446 -198 447 -197
rect 447 -198 448 -197
rect 448 -198 449 -197
rect 449 -198 450 -197
rect 450 -198 451 -197
rect 451 -198 452 -197
rect 452 -198 453 -197
rect 453 -198 454 -197
rect 454 -198 455 -197
rect 455 -198 456 -197
rect 456 -198 457 -197
rect 457 -198 458 -197
rect 458 -198 459 -197
rect 459 -198 460 -197
rect 460 -198 461 -197
rect 461 -198 462 -197
rect 462 -198 463 -197
rect 463 -198 464 -197
rect 464 -198 465 -197
rect 465 -198 466 -197
rect 466 -198 467 -197
rect 467 -198 468 -197
rect 468 -198 469 -197
rect 469 -198 470 -197
rect 470 -198 471 -197
rect 471 -198 472 -197
rect 472 -198 473 -197
rect 473 -198 474 -197
rect 474 -198 475 -197
rect 475 -198 476 -197
rect 476 -198 477 -197
rect 477 -198 478 -197
rect 478 -198 479 -197
rect 479 -198 480 -197
rect 2 -199 3 -198
rect 3 -199 4 -198
rect 4 -199 5 -198
rect 5 -199 6 -198
rect 6 -199 7 -198
rect 7 -199 8 -198
rect 8 -199 9 -198
rect 9 -199 10 -198
rect 10 -199 11 -198
rect 11 -199 12 -198
rect 12 -199 13 -198
rect 13 -199 14 -198
rect 14 -199 15 -198
rect 15 -199 16 -198
rect 16 -199 17 -198
rect 17 -199 18 -198
rect 18 -199 19 -198
rect 19 -199 20 -198
rect 20 -199 21 -198
rect 21 -199 22 -198
rect 22 -199 23 -198
rect 23 -199 24 -198
rect 24 -199 25 -198
rect 25 -199 26 -198
rect 26 -199 27 -198
rect 27 -199 28 -198
rect 28 -199 29 -198
rect 29 -199 30 -198
rect 30 -199 31 -198
rect 31 -199 32 -198
rect 32 -199 33 -198
rect 33 -199 34 -198
rect 34 -199 35 -198
rect 35 -199 36 -198
rect 36 -199 37 -198
rect 37 -199 38 -198
rect 38 -199 39 -198
rect 39 -199 40 -198
rect 40 -199 41 -198
rect 41 -199 42 -198
rect 42 -199 43 -198
rect 43 -199 44 -198
rect 44 -199 45 -198
rect 45 -199 46 -198
rect 46 -199 47 -198
rect 47 -199 48 -198
rect 48 -199 49 -198
rect 49 -199 50 -198
rect 50 -199 51 -198
rect 51 -199 52 -198
rect 52 -199 53 -198
rect 53 -199 54 -198
rect 54 -199 55 -198
rect 55 -199 56 -198
rect 56 -199 57 -198
rect 57 -199 58 -198
rect 58 -199 59 -198
rect 59 -199 60 -198
rect 60 -199 61 -198
rect 61 -199 62 -198
rect 62 -199 63 -198
rect 63 -199 64 -198
rect 64 -199 65 -198
rect 65 -199 66 -198
rect 66 -199 67 -198
rect 67 -199 68 -198
rect 68 -199 69 -198
rect 69 -199 70 -198
rect 70 -199 71 -198
rect 71 -199 72 -198
rect 72 -199 73 -198
rect 73 -199 74 -198
rect 74 -199 75 -198
rect 75 -199 76 -198
rect 76 -199 77 -198
rect 77 -199 78 -198
rect 78 -199 79 -198
rect 79 -199 80 -198
rect 80 -199 81 -198
rect 81 -199 82 -198
rect 82 -199 83 -198
rect 83 -199 84 -198
rect 84 -199 85 -198
rect 85 -199 86 -198
rect 86 -199 87 -198
rect 87 -199 88 -198
rect 88 -199 89 -198
rect 89 -199 90 -198
rect 90 -199 91 -198
rect 91 -199 92 -198
rect 92 -199 93 -198
rect 93 -199 94 -198
rect 94 -199 95 -198
rect 95 -199 96 -198
rect 96 -199 97 -198
rect 97 -199 98 -198
rect 98 -199 99 -198
rect 99 -199 100 -198
rect 100 -199 101 -198
rect 101 -199 102 -198
rect 102 -199 103 -198
rect 103 -199 104 -198
rect 104 -199 105 -198
rect 105 -199 106 -198
rect 106 -199 107 -198
rect 107 -199 108 -198
rect 108 -199 109 -198
rect 109 -199 110 -198
rect 110 -199 111 -198
rect 111 -199 112 -198
rect 112 -199 113 -198
rect 113 -199 114 -198
rect 114 -199 115 -198
rect 115 -199 116 -198
rect 116 -199 117 -198
rect 117 -199 118 -198
rect 118 -199 119 -198
rect 119 -199 120 -198
rect 120 -199 121 -198
rect 121 -199 122 -198
rect 122 -199 123 -198
rect 123 -199 124 -198
rect 124 -199 125 -198
rect 125 -199 126 -198
rect 126 -199 127 -198
rect 127 -199 128 -198
rect 128 -199 129 -198
rect 129 -199 130 -198
rect 130 -199 131 -198
rect 131 -199 132 -198
rect 132 -199 133 -198
rect 133 -199 134 -198
rect 134 -199 135 -198
rect 135 -199 136 -198
rect 136 -199 137 -198
rect 137 -199 138 -198
rect 138 -199 139 -198
rect 139 -199 140 -198
rect 140 -199 141 -198
rect 141 -199 142 -198
rect 142 -199 143 -198
rect 143 -199 144 -198
rect 144 -199 145 -198
rect 145 -199 146 -198
rect 146 -199 147 -198
rect 147 -199 148 -198
rect 148 -199 149 -198
rect 149 -199 150 -198
rect 150 -199 151 -198
rect 151 -199 152 -198
rect 152 -199 153 -198
rect 153 -199 154 -198
rect 154 -199 155 -198
rect 155 -199 156 -198
rect 156 -199 157 -198
rect 157 -199 158 -198
rect 158 -199 159 -198
rect 159 -199 160 -198
rect 160 -199 161 -198
rect 161 -199 162 -198
rect 162 -199 163 -198
rect 163 -199 164 -198
rect 164 -199 165 -198
rect 165 -199 166 -198
rect 166 -199 167 -198
rect 167 -199 168 -198
rect 168 -199 169 -198
rect 169 -199 170 -198
rect 170 -199 171 -198
rect 171 -199 172 -198
rect 172 -199 173 -198
rect 173 -199 174 -198
rect 174 -199 175 -198
rect 175 -199 176 -198
rect 176 -199 177 -198
rect 177 -199 178 -198
rect 178 -199 179 -198
rect 179 -199 180 -198
rect 180 -199 181 -198
rect 181 -199 182 -198
rect 182 -199 183 -198
rect 183 -199 184 -198
rect 184 -199 185 -198
rect 185 -199 186 -198
rect 186 -199 187 -198
rect 187 -199 188 -198
rect 188 -199 189 -198
rect 189 -199 190 -198
rect 190 -199 191 -198
rect 191 -199 192 -198
rect 192 -199 193 -198
rect 193 -199 194 -198
rect 194 -199 195 -198
rect 195 -199 196 -198
rect 196 -199 197 -198
rect 197 -199 198 -198
rect 198 -199 199 -198
rect 199 -199 200 -198
rect 200 -199 201 -198
rect 201 -199 202 -198
rect 202 -199 203 -198
rect 203 -199 204 -198
rect 204 -199 205 -198
rect 205 -199 206 -198
rect 206 -199 207 -198
rect 207 -199 208 -198
rect 208 -199 209 -198
rect 209 -199 210 -198
rect 210 -199 211 -198
rect 211 -199 212 -198
rect 212 -199 213 -198
rect 213 -199 214 -198
rect 214 -199 215 -198
rect 215 -199 216 -198
rect 216 -199 217 -198
rect 217 -199 218 -198
rect 218 -199 219 -198
rect 219 -199 220 -198
rect 220 -199 221 -198
rect 221 -199 222 -198
rect 222 -199 223 -198
rect 223 -199 224 -198
rect 224 -199 225 -198
rect 225 -199 226 -198
rect 226 -199 227 -198
rect 227 -199 228 -198
rect 228 -199 229 -198
rect 229 -199 230 -198
rect 230 -199 231 -198
rect 231 -199 232 -198
rect 232 -199 233 -198
rect 233 -199 234 -198
rect 234 -199 235 -198
rect 235 -199 236 -198
rect 236 -199 237 -198
rect 237 -199 238 -198
rect 238 -199 239 -198
rect 239 -199 240 -198
rect 240 -199 241 -198
rect 241 -199 242 -198
rect 242 -199 243 -198
rect 243 -199 244 -198
rect 244 -199 245 -198
rect 245 -199 246 -198
rect 246 -199 247 -198
rect 247 -199 248 -198
rect 248 -199 249 -198
rect 249 -199 250 -198
rect 250 -199 251 -198
rect 251 -199 252 -198
rect 252 -199 253 -198
rect 253 -199 254 -198
rect 254 -199 255 -198
rect 255 -199 256 -198
rect 256 -199 257 -198
rect 257 -199 258 -198
rect 258 -199 259 -198
rect 259 -199 260 -198
rect 260 -199 261 -198
rect 261 -199 262 -198
rect 262 -199 263 -198
rect 263 -199 264 -198
rect 264 -199 265 -198
rect 265 -199 266 -198
rect 266 -199 267 -198
rect 267 -199 268 -198
rect 268 -199 269 -198
rect 269 -199 270 -198
rect 270 -199 271 -198
rect 271 -199 272 -198
rect 272 -199 273 -198
rect 273 -199 274 -198
rect 274 -199 275 -198
rect 275 -199 276 -198
rect 276 -199 277 -198
rect 277 -199 278 -198
rect 278 -199 279 -198
rect 279 -199 280 -198
rect 280 -199 281 -198
rect 281 -199 282 -198
rect 282 -199 283 -198
rect 283 -199 284 -198
rect 284 -199 285 -198
rect 285 -199 286 -198
rect 286 -199 287 -198
rect 287 -199 288 -198
rect 288 -199 289 -198
rect 289 -199 290 -198
rect 290 -199 291 -198
rect 291 -199 292 -198
rect 292 -199 293 -198
rect 293 -199 294 -198
rect 294 -199 295 -198
rect 295 -199 296 -198
rect 296 -199 297 -198
rect 297 -199 298 -198
rect 298 -199 299 -198
rect 299 -199 300 -198
rect 300 -199 301 -198
rect 301 -199 302 -198
rect 302 -199 303 -198
rect 303 -199 304 -198
rect 304 -199 305 -198
rect 305 -199 306 -198
rect 306 -199 307 -198
rect 307 -199 308 -198
rect 308 -199 309 -198
rect 309 -199 310 -198
rect 310 -199 311 -198
rect 311 -199 312 -198
rect 312 -199 313 -198
rect 313 -199 314 -198
rect 314 -199 315 -198
rect 315 -199 316 -198
rect 316 -199 317 -198
rect 317 -199 318 -198
rect 318 -199 319 -198
rect 319 -199 320 -198
rect 320 -199 321 -198
rect 321 -199 322 -198
rect 322 -199 323 -198
rect 323 -199 324 -198
rect 324 -199 325 -198
rect 325 -199 326 -198
rect 326 -199 327 -198
rect 327 -199 328 -198
rect 328 -199 329 -198
rect 329 -199 330 -198
rect 330 -199 331 -198
rect 331 -199 332 -198
rect 332 -199 333 -198
rect 333 -199 334 -198
rect 334 -199 335 -198
rect 335 -199 336 -198
rect 336 -199 337 -198
rect 337 -199 338 -198
rect 338 -199 339 -198
rect 339 -199 340 -198
rect 340 -199 341 -198
rect 341 -199 342 -198
rect 342 -199 343 -198
rect 343 -199 344 -198
rect 344 -199 345 -198
rect 345 -199 346 -198
rect 346 -199 347 -198
rect 347 -199 348 -198
rect 348 -199 349 -198
rect 349 -199 350 -198
rect 350 -199 351 -198
rect 351 -199 352 -198
rect 352 -199 353 -198
rect 353 -199 354 -198
rect 354 -199 355 -198
rect 355 -199 356 -198
rect 356 -199 357 -198
rect 357 -199 358 -198
rect 358 -199 359 -198
rect 359 -199 360 -198
rect 360 -199 361 -198
rect 361 -199 362 -198
rect 362 -199 363 -198
rect 363 -199 364 -198
rect 364 -199 365 -198
rect 365 -199 366 -198
rect 366 -199 367 -198
rect 367 -199 368 -198
rect 368 -199 369 -198
rect 369 -199 370 -198
rect 370 -199 371 -198
rect 371 -199 372 -198
rect 372 -199 373 -198
rect 373 -199 374 -198
rect 374 -199 375 -198
rect 375 -199 376 -198
rect 376 -199 377 -198
rect 377 -199 378 -198
rect 378 -199 379 -198
rect 379 -199 380 -198
rect 380 -199 381 -198
rect 381 -199 382 -198
rect 382 -199 383 -198
rect 383 -199 384 -198
rect 384 -199 385 -198
rect 385 -199 386 -198
rect 386 -199 387 -198
rect 387 -199 388 -198
rect 388 -199 389 -198
rect 389 -199 390 -198
rect 390 -199 391 -198
rect 391 -199 392 -198
rect 392 -199 393 -198
rect 393 -199 394 -198
rect 394 -199 395 -198
rect 395 -199 396 -198
rect 396 -199 397 -198
rect 397 -199 398 -198
rect 398 -199 399 -198
rect 399 -199 400 -198
rect 400 -199 401 -198
rect 401 -199 402 -198
rect 402 -199 403 -198
rect 403 -199 404 -198
rect 404 -199 405 -198
rect 405 -199 406 -198
rect 406 -199 407 -198
rect 407 -199 408 -198
rect 408 -199 409 -198
rect 409 -199 410 -198
rect 410 -199 411 -198
rect 411 -199 412 -198
rect 412 -199 413 -198
rect 413 -199 414 -198
rect 414 -199 415 -198
rect 415 -199 416 -198
rect 416 -199 417 -198
rect 417 -199 418 -198
rect 418 -199 419 -198
rect 419 -199 420 -198
rect 420 -199 421 -198
rect 421 -199 422 -198
rect 422 -199 423 -198
rect 423 -199 424 -198
rect 424 -199 425 -198
rect 425 -199 426 -198
rect 426 -199 427 -198
rect 427 -199 428 -198
rect 428 -199 429 -198
rect 429 -199 430 -198
rect 430 -199 431 -198
rect 431 -199 432 -198
rect 432 -199 433 -198
rect 433 -199 434 -198
rect 434 -199 435 -198
rect 435 -199 436 -198
rect 436 -199 437 -198
rect 437 -199 438 -198
rect 438 -199 439 -198
rect 439 -199 440 -198
rect 440 -199 441 -198
rect 441 -199 442 -198
rect 442 -199 443 -198
rect 443 -199 444 -198
rect 444 -199 445 -198
rect 445 -199 446 -198
rect 446 -199 447 -198
rect 447 -199 448 -198
rect 448 -199 449 -198
rect 449 -199 450 -198
rect 450 -199 451 -198
rect 451 -199 452 -198
rect 452 -199 453 -198
rect 453 -199 454 -198
rect 454 -199 455 -198
rect 455 -199 456 -198
rect 456 -199 457 -198
rect 457 -199 458 -198
rect 458 -199 459 -198
rect 459 -199 460 -198
rect 460 -199 461 -198
rect 461 -199 462 -198
rect 462 -199 463 -198
rect 463 -199 464 -198
rect 464 -199 465 -198
rect 465 -199 466 -198
rect 466 -199 467 -198
rect 467 -199 468 -198
rect 468 -199 469 -198
rect 469 -199 470 -198
rect 470 -199 471 -198
rect 471 -199 472 -198
rect 472 -199 473 -198
rect 473 -199 474 -198
rect 474 -199 475 -198
rect 475 -199 476 -198
rect 476 -199 477 -198
rect 477 -199 478 -198
rect 478 -199 479 -198
rect 479 -199 480 -198
rect 2 -200 3 -199
rect 3 -200 4 -199
rect 4 -200 5 -199
rect 5 -200 6 -199
rect 6 -200 7 -199
rect 7 -200 8 -199
rect 8 -200 9 -199
rect 9 -200 10 -199
rect 10 -200 11 -199
rect 11 -200 12 -199
rect 12 -200 13 -199
rect 13 -200 14 -199
rect 14 -200 15 -199
rect 15 -200 16 -199
rect 16 -200 17 -199
rect 17 -200 18 -199
rect 18 -200 19 -199
rect 19 -200 20 -199
rect 20 -200 21 -199
rect 21 -200 22 -199
rect 22 -200 23 -199
rect 23 -200 24 -199
rect 24 -200 25 -199
rect 25 -200 26 -199
rect 26 -200 27 -199
rect 27 -200 28 -199
rect 28 -200 29 -199
rect 29 -200 30 -199
rect 30 -200 31 -199
rect 31 -200 32 -199
rect 32 -200 33 -199
rect 33 -200 34 -199
rect 34 -200 35 -199
rect 35 -200 36 -199
rect 36 -200 37 -199
rect 37 -200 38 -199
rect 38 -200 39 -199
rect 39 -200 40 -199
rect 40 -200 41 -199
rect 41 -200 42 -199
rect 42 -200 43 -199
rect 43 -200 44 -199
rect 44 -200 45 -199
rect 45 -200 46 -199
rect 46 -200 47 -199
rect 47 -200 48 -199
rect 48 -200 49 -199
rect 49 -200 50 -199
rect 50 -200 51 -199
rect 51 -200 52 -199
rect 52 -200 53 -199
rect 53 -200 54 -199
rect 54 -200 55 -199
rect 55 -200 56 -199
rect 56 -200 57 -199
rect 57 -200 58 -199
rect 58 -200 59 -199
rect 59 -200 60 -199
rect 60 -200 61 -199
rect 61 -200 62 -199
rect 62 -200 63 -199
rect 63 -200 64 -199
rect 64 -200 65 -199
rect 65 -200 66 -199
rect 66 -200 67 -199
rect 67 -200 68 -199
rect 68 -200 69 -199
rect 69 -200 70 -199
rect 70 -200 71 -199
rect 71 -200 72 -199
rect 72 -200 73 -199
rect 73 -200 74 -199
rect 74 -200 75 -199
rect 75 -200 76 -199
rect 76 -200 77 -199
rect 77 -200 78 -199
rect 78 -200 79 -199
rect 79 -200 80 -199
rect 80 -200 81 -199
rect 81 -200 82 -199
rect 82 -200 83 -199
rect 83 -200 84 -199
rect 84 -200 85 -199
rect 85 -200 86 -199
rect 86 -200 87 -199
rect 87 -200 88 -199
rect 88 -200 89 -199
rect 89 -200 90 -199
rect 90 -200 91 -199
rect 91 -200 92 -199
rect 92 -200 93 -199
rect 93 -200 94 -199
rect 94 -200 95 -199
rect 95 -200 96 -199
rect 96 -200 97 -199
rect 97 -200 98 -199
rect 98 -200 99 -199
rect 99 -200 100 -199
rect 100 -200 101 -199
rect 101 -200 102 -199
rect 102 -200 103 -199
rect 103 -200 104 -199
rect 104 -200 105 -199
rect 105 -200 106 -199
rect 106 -200 107 -199
rect 107 -200 108 -199
rect 108 -200 109 -199
rect 109 -200 110 -199
rect 110 -200 111 -199
rect 111 -200 112 -199
rect 112 -200 113 -199
rect 113 -200 114 -199
rect 114 -200 115 -199
rect 115 -200 116 -199
rect 116 -200 117 -199
rect 117 -200 118 -199
rect 118 -200 119 -199
rect 119 -200 120 -199
rect 120 -200 121 -199
rect 121 -200 122 -199
rect 122 -200 123 -199
rect 123 -200 124 -199
rect 124 -200 125 -199
rect 125 -200 126 -199
rect 126 -200 127 -199
rect 127 -200 128 -199
rect 128 -200 129 -199
rect 129 -200 130 -199
rect 130 -200 131 -199
rect 131 -200 132 -199
rect 132 -200 133 -199
rect 133 -200 134 -199
rect 134 -200 135 -199
rect 135 -200 136 -199
rect 136 -200 137 -199
rect 137 -200 138 -199
rect 138 -200 139 -199
rect 139 -200 140 -199
rect 140 -200 141 -199
rect 141 -200 142 -199
rect 142 -200 143 -199
rect 143 -200 144 -199
rect 144 -200 145 -199
rect 145 -200 146 -199
rect 146 -200 147 -199
rect 147 -200 148 -199
rect 148 -200 149 -199
rect 149 -200 150 -199
rect 150 -200 151 -199
rect 151 -200 152 -199
rect 152 -200 153 -199
rect 153 -200 154 -199
rect 154 -200 155 -199
rect 155 -200 156 -199
rect 156 -200 157 -199
rect 157 -200 158 -199
rect 158 -200 159 -199
rect 159 -200 160 -199
rect 160 -200 161 -199
rect 161 -200 162 -199
rect 162 -200 163 -199
rect 163 -200 164 -199
rect 164 -200 165 -199
rect 165 -200 166 -199
rect 166 -200 167 -199
rect 167 -200 168 -199
rect 168 -200 169 -199
rect 169 -200 170 -199
rect 170 -200 171 -199
rect 171 -200 172 -199
rect 172 -200 173 -199
rect 173 -200 174 -199
rect 174 -200 175 -199
rect 175 -200 176 -199
rect 176 -200 177 -199
rect 177 -200 178 -199
rect 178 -200 179 -199
rect 179 -200 180 -199
rect 180 -200 181 -199
rect 181 -200 182 -199
rect 182 -200 183 -199
rect 183 -200 184 -199
rect 184 -200 185 -199
rect 185 -200 186 -199
rect 186 -200 187 -199
rect 187 -200 188 -199
rect 188 -200 189 -199
rect 189 -200 190 -199
rect 190 -200 191 -199
rect 191 -200 192 -199
rect 192 -200 193 -199
rect 193 -200 194 -199
rect 194 -200 195 -199
rect 195 -200 196 -199
rect 196 -200 197 -199
rect 197 -200 198 -199
rect 198 -200 199 -199
rect 199 -200 200 -199
rect 200 -200 201 -199
rect 201 -200 202 -199
rect 202 -200 203 -199
rect 203 -200 204 -199
rect 204 -200 205 -199
rect 205 -200 206 -199
rect 206 -200 207 -199
rect 207 -200 208 -199
rect 208 -200 209 -199
rect 209 -200 210 -199
rect 210 -200 211 -199
rect 211 -200 212 -199
rect 212 -200 213 -199
rect 213 -200 214 -199
rect 214 -200 215 -199
rect 215 -200 216 -199
rect 216 -200 217 -199
rect 217 -200 218 -199
rect 218 -200 219 -199
rect 219 -200 220 -199
rect 220 -200 221 -199
rect 221 -200 222 -199
rect 222 -200 223 -199
rect 223 -200 224 -199
rect 224 -200 225 -199
rect 225 -200 226 -199
rect 226 -200 227 -199
rect 227 -200 228 -199
rect 228 -200 229 -199
rect 229 -200 230 -199
rect 230 -200 231 -199
rect 231 -200 232 -199
rect 232 -200 233 -199
rect 233 -200 234 -199
rect 234 -200 235 -199
rect 235 -200 236 -199
rect 236 -200 237 -199
rect 237 -200 238 -199
rect 238 -200 239 -199
rect 239 -200 240 -199
rect 240 -200 241 -199
rect 241 -200 242 -199
rect 242 -200 243 -199
rect 243 -200 244 -199
rect 244 -200 245 -199
rect 245 -200 246 -199
rect 246 -200 247 -199
rect 247 -200 248 -199
rect 248 -200 249 -199
rect 249 -200 250 -199
rect 250 -200 251 -199
rect 251 -200 252 -199
rect 252 -200 253 -199
rect 253 -200 254 -199
rect 254 -200 255 -199
rect 255 -200 256 -199
rect 256 -200 257 -199
rect 257 -200 258 -199
rect 258 -200 259 -199
rect 259 -200 260 -199
rect 260 -200 261 -199
rect 261 -200 262 -199
rect 262 -200 263 -199
rect 263 -200 264 -199
rect 264 -200 265 -199
rect 265 -200 266 -199
rect 266 -200 267 -199
rect 267 -200 268 -199
rect 268 -200 269 -199
rect 269 -200 270 -199
rect 270 -200 271 -199
rect 271 -200 272 -199
rect 272 -200 273 -199
rect 273 -200 274 -199
rect 274 -200 275 -199
rect 275 -200 276 -199
rect 276 -200 277 -199
rect 277 -200 278 -199
rect 278 -200 279 -199
rect 279 -200 280 -199
rect 280 -200 281 -199
rect 281 -200 282 -199
rect 282 -200 283 -199
rect 283 -200 284 -199
rect 284 -200 285 -199
rect 285 -200 286 -199
rect 286 -200 287 -199
rect 287 -200 288 -199
rect 288 -200 289 -199
rect 289 -200 290 -199
rect 290 -200 291 -199
rect 291 -200 292 -199
rect 292 -200 293 -199
rect 293 -200 294 -199
rect 294 -200 295 -199
rect 295 -200 296 -199
rect 296 -200 297 -199
rect 297 -200 298 -199
rect 298 -200 299 -199
rect 299 -200 300 -199
rect 300 -200 301 -199
rect 301 -200 302 -199
rect 302 -200 303 -199
rect 303 -200 304 -199
rect 304 -200 305 -199
rect 305 -200 306 -199
rect 306 -200 307 -199
rect 307 -200 308 -199
rect 308 -200 309 -199
rect 309 -200 310 -199
rect 310 -200 311 -199
rect 311 -200 312 -199
rect 312 -200 313 -199
rect 313 -200 314 -199
rect 314 -200 315 -199
rect 315 -200 316 -199
rect 316 -200 317 -199
rect 317 -200 318 -199
rect 318 -200 319 -199
rect 319 -200 320 -199
rect 320 -200 321 -199
rect 321 -200 322 -199
rect 322 -200 323 -199
rect 323 -200 324 -199
rect 324 -200 325 -199
rect 325 -200 326 -199
rect 326 -200 327 -199
rect 327 -200 328 -199
rect 328 -200 329 -199
rect 329 -200 330 -199
rect 330 -200 331 -199
rect 331 -200 332 -199
rect 332 -200 333 -199
rect 333 -200 334 -199
rect 334 -200 335 -199
rect 335 -200 336 -199
rect 336 -200 337 -199
rect 337 -200 338 -199
rect 338 -200 339 -199
rect 339 -200 340 -199
rect 340 -200 341 -199
rect 341 -200 342 -199
rect 342 -200 343 -199
rect 343 -200 344 -199
rect 344 -200 345 -199
rect 345 -200 346 -199
rect 346 -200 347 -199
rect 347 -200 348 -199
rect 348 -200 349 -199
rect 349 -200 350 -199
rect 350 -200 351 -199
rect 351 -200 352 -199
rect 352 -200 353 -199
rect 353 -200 354 -199
rect 354 -200 355 -199
rect 355 -200 356 -199
rect 356 -200 357 -199
rect 357 -200 358 -199
rect 358 -200 359 -199
rect 359 -200 360 -199
rect 360 -200 361 -199
rect 361 -200 362 -199
rect 362 -200 363 -199
rect 363 -200 364 -199
rect 364 -200 365 -199
rect 365 -200 366 -199
rect 366 -200 367 -199
rect 367 -200 368 -199
rect 368 -200 369 -199
rect 369 -200 370 -199
rect 370 -200 371 -199
rect 371 -200 372 -199
rect 372 -200 373 -199
rect 373 -200 374 -199
rect 374 -200 375 -199
rect 375 -200 376 -199
rect 376 -200 377 -199
rect 377 -200 378 -199
rect 378 -200 379 -199
rect 379 -200 380 -199
rect 380 -200 381 -199
rect 381 -200 382 -199
rect 382 -200 383 -199
rect 383 -200 384 -199
rect 384 -200 385 -199
rect 385 -200 386 -199
rect 386 -200 387 -199
rect 387 -200 388 -199
rect 388 -200 389 -199
rect 389 -200 390 -199
rect 390 -200 391 -199
rect 391 -200 392 -199
rect 392 -200 393 -199
rect 393 -200 394 -199
rect 394 -200 395 -199
rect 395 -200 396 -199
rect 396 -200 397 -199
rect 397 -200 398 -199
rect 398 -200 399 -199
rect 399 -200 400 -199
rect 400 -200 401 -199
rect 401 -200 402 -199
rect 402 -200 403 -199
rect 403 -200 404 -199
rect 404 -200 405 -199
rect 405 -200 406 -199
rect 406 -200 407 -199
rect 407 -200 408 -199
rect 408 -200 409 -199
rect 409 -200 410 -199
rect 410 -200 411 -199
rect 411 -200 412 -199
rect 412 -200 413 -199
rect 413 -200 414 -199
rect 414 -200 415 -199
rect 415 -200 416 -199
rect 416 -200 417 -199
rect 417 -200 418 -199
rect 418 -200 419 -199
rect 419 -200 420 -199
rect 420 -200 421 -199
rect 421 -200 422 -199
rect 422 -200 423 -199
rect 423 -200 424 -199
rect 424 -200 425 -199
rect 425 -200 426 -199
rect 426 -200 427 -199
rect 427 -200 428 -199
rect 428 -200 429 -199
rect 429 -200 430 -199
rect 430 -200 431 -199
rect 431 -200 432 -199
rect 432 -200 433 -199
rect 433 -200 434 -199
rect 434 -200 435 -199
rect 435 -200 436 -199
rect 436 -200 437 -199
rect 437 -200 438 -199
rect 438 -200 439 -199
rect 439 -200 440 -199
rect 440 -200 441 -199
rect 441 -200 442 -199
rect 442 -200 443 -199
rect 443 -200 444 -199
rect 444 -200 445 -199
rect 445 -200 446 -199
rect 446 -200 447 -199
rect 447 -200 448 -199
rect 448 -200 449 -199
rect 449 -200 450 -199
rect 450 -200 451 -199
rect 451 -200 452 -199
rect 452 -200 453 -199
rect 453 -200 454 -199
rect 454 -200 455 -199
rect 455 -200 456 -199
rect 456 -200 457 -199
rect 457 -200 458 -199
rect 458 -200 459 -199
rect 459 -200 460 -199
rect 460 -200 461 -199
rect 461 -200 462 -199
rect 462 -200 463 -199
rect 463 -200 464 -199
rect 464 -200 465 -199
rect 465 -200 466 -199
rect 466 -200 467 -199
rect 467 -200 468 -199
rect 468 -200 469 -199
rect 469 -200 470 -199
rect 470 -200 471 -199
rect 471 -200 472 -199
rect 472 -200 473 -199
rect 473 -200 474 -199
rect 474 -200 475 -199
rect 475 -200 476 -199
rect 476 -200 477 -199
rect 477 -200 478 -199
rect 478 -200 479 -199
rect 479 -200 480 -199
rect 2 -201 3 -200
rect 3 -201 4 -200
rect 4 -201 5 -200
rect 5 -201 6 -200
rect 6 -201 7 -200
rect 7 -201 8 -200
rect 8 -201 9 -200
rect 9 -201 10 -200
rect 10 -201 11 -200
rect 11 -201 12 -200
rect 12 -201 13 -200
rect 13 -201 14 -200
rect 14 -201 15 -200
rect 15 -201 16 -200
rect 16 -201 17 -200
rect 17 -201 18 -200
rect 18 -201 19 -200
rect 19 -201 20 -200
rect 20 -201 21 -200
rect 21 -201 22 -200
rect 22 -201 23 -200
rect 23 -201 24 -200
rect 24 -201 25 -200
rect 25 -201 26 -200
rect 26 -201 27 -200
rect 27 -201 28 -200
rect 28 -201 29 -200
rect 29 -201 30 -200
rect 30 -201 31 -200
rect 31 -201 32 -200
rect 32 -201 33 -200
rect 33 -201 34 -200
rect 34 -201 35 -200
rect 35 -201 36 -200
rect 36 -201 37 -200
rect 37 -201 38 -200
rect 38 -201 39 -200
rect 39 -201 40 -200
rect 40 -201 41 -200
rect 41 -201 42 -200
rect 42 -201 43 -200
rect 43 -201 44 -200
rect 44 -201 45 -200
rect 45 -201 46 -200
rect 46 -201 47 -200
rect 47 -201 48 -200
rect 48 -201 49 -200
rect 49 -201 50 -200
rect 50 -201 51 -200
rect 51 -201 52 -200
rect 52 -201 53 -200
rect 53 -201 54 -200
rect 54 -201 55 -200
rect 55 -201 56 -200
rect 56 -201 57 -200
rect 57 -201 58 -200
rect 58 -201 59 -200
rect 59 -201 60 -200
rect 60 -201 61 -200
rect 61 -201 62 -200
rect 62 -201 63 -200
rect 63 -201 64 -200
rect 64 -201 65 -200
rect 65 -201 66 -200
rect 66 -201 67 -200
rect 67 -201 68 -200
rect 68 -201 69 -200
rect 69 -201 70 -200
rect 70 -201 71 -200
rect 71 -201 72 -200
rect 72 -201 73 -200
rect 73 -201 74 -200
rect 74 -201 75 -200
rect 75 -201 76 -200
rect 76 -201 77 -200
rect 77 -201 78 -200
rect 78 -201 79 -200
rect 79 -201 80 -200
rect 80 -201 81 -200
rect 81 -201 82 -200
rect 82 -201 83 -200
rect 83 -201 84 -200
rect 84 -201 85 -200
rect 85 -201 86 -200
rect 86 -201 87 -200
rect 87 -201 88 -200
rect 88 -201 89 -200
rect 89 -201 90 -200
rect 90 -201 91 -200
rect 91 -201 92 -200
rect 92 -201 93 -200
rect 93 -201 94 -200
rect 94 -201 95 -200
rect 95 -201 96 -200
rect 96 -201 97 -200
rect 97 -201 98 -200
rect 98 -201 99 -200
rect 99 -201 100 -200
rect 100 -201 101 -200
rect 101 -201 102 -200
rect 102 -201 103 -200
rect 103 -201 104 -200
rect 104 -201 105 -200
rect 105 -201 106 -200
rect 106 -201 107 -200
rect 107 -201 108 -200
rect 108 -201 109 -200
rect 109 -201 110 -200
rect 110 -201 111 -200
rect 111 -201 112 -200
rect 112 -201 113 -200
rect 113 -201 114 -200
rect 114 -201 115 -200
rect 115 -201 116 -200
rect 116 -201 117 -200
rect 117 -201 118 -200
rect 118 -201 119 -200
rect 119 -201 120 -200
rect 120 -201 121 -200
rect 121 -201 122 -200
rect 122 -201 123 -200
rect 123 -201 124 -200
rect 124 -201 125 -200
rect 125 -201 126 -200
rect 126 -201 127 -200
rect 127 -201 128 -200
rect 128 -201 129 -200
rect 129 -201 130 -200
rect 130 -201 131 -200
rect 131 -201 132 -200
rect 132 -201 133 -200
rect 133 -201 134 -200
rect 134 -201 135 -200
rect 135 -201 136 -200
rect 136 -201 137 -200
rect 137 -201 138 -200
rect 138 -201 139 -200
rect 139 -201 140 -200
rect 140 -201 141 -200
rect 141 -201 142 -200
rect 142 -201 143 -200
rect 143 -201 144 -200
rect 144 -201 145 -200
rect 145 -201 146 -200
rect 146 -201 147 -200
rect 147 -201 148 -200
rect 148 -201 149 -200
rect 149 -201 150 -200
rect 150 -201 151 -200
rect 151 -201 152 -200
rect 152 -201 153 -200
rect 153 -201 154 -200
rect 154 -201 155 -200
rect 155 -201 156 -200
rect 156 -201 157 -200
rect 157 -201 158 -200
rect 158 -201 159 -200
rect 159 -201 160 -200
rect 160 -201 161 -200
rect 161 -201 162 -200
rect 162 -201 163 -200
rect 163 -201 164 -200
rect 164 -201 165 -200
rect 165 -201 166 -200
rect 166 -201 167 -200
rect 167 -201 168 -200
rect 168 -201 169 -200
rect 169 -201 170 -200
rect 170 -201 171 -200
rect 171 -201 172 -200
rect 172 -201 173 -200
rect 173 -201 174 -200
rect 174 -201 175 -200
rect 175 -201 176 -200
rect 176 -201 177 -200
rect 177 -201 178 -200
rect 178 -201 179 -200
rect 179 -201 180 -200
rect 180 -201 181 -200
rect 181 -201 182 -200
rect 182 -201 183 -200
rect 183 -201 184 -200
rect 184 -201 185 -200
rect 185 -201 186 -200
rect 186 -201 187 -200
rect 187 -201 188 -200
rect 188 -201 189 -200
rect 189 -201 190 -200
rect 190 -201 191 -200
rect 191 -201 192 -200
rect 192 -201 193 -200
rect 193 -201 194 -200
rect 194 -201 195 -200
rect 195 -201 196 -200
rect 196 -201 197 -200
rect 197 -201 198 -200
rect 198 -201 199 -200
rect 199 -201 200 -200
rect 200 -201 201 -200
rect 201 -201 202 -200
rect 202 -201 203 -200
rect 203 -201 204 -200
rect 204 -201 205 -200
rect 205 -201 206 -200
rect 206 -201 207 -200
rect 207 -201 208 -200
rect 208 -201 209 -200
rect 209 -201 210 -200
rect 210 -201 211 -200
rect 211 -201 212 -200
rect 212 -201 213 -200
rect 213 -201 214 -200
rect 214 -201 215 -200
rect 215 -201 216 -200
rect 216 -201 217 -200
rect 217 -201 218 -200
rect 218 -201 219 -200
rect 219 -201 220 -200
rect 220 -201 221 -200
rect 221 -201 222 -200
rect 222 -201 223 -200
rect 223 -201 224 -200
rect 224 -201 225 -200
rect 225 -201 226 -200
rect 226 -201 227 -200
rect 227 -201 228 -200
rect 228 -201 229 -200
rect 229 -201 230 -200
rect 230 -201 231 -200
rect 231 -201 232 -200
rect 232 -201 233 -200
rect 233 -201 234 -200
rect 234 -201 235 -200
rect 235 -201 236 -200
rect 236 -201 237 -200
rect 237 -201 238 -200
rect 238 -201 239 -200
rect 239 -201 240 -200
rect 240 -201 241 -200
rect 241 -201 242 -200
rect 242 -201 243 -200
rect 243 -201 244 -200
rect 244 -201 245 -200
rect 245 -201 246 -200
rect 246 -201 247 -200
rect 247 -201 248 -200
rect 248 -201 249 -200
rect 249 -201 250 -200
rect 250 -201 251 -200
rect 251 -201 252 -200
rect 252 -201 253 -200
rect 253 -201 254 -200
rect 254 -201 255 -200
rect 255 -201 256 -200
rect 256 -201 257 -200
rect 257 -201 258 -200
rect 258 -201 259 -200
rect 259 -201 260 -200
rect 260 -201 261 -200
rect 261 -201 262 -200
rect 262 -201 263 -200
rect 263 -201 264 -200
rect 264 -201 265 -200
rect 265 -201 266 -200
rect 266 -201 267 -200
rect 267 -201 268 -200
rect 268 -201 269 -200
rect 269 -201 270 -200
rect 270 -201 271 -200
rect 271 -201 272 -200
rect 272 -201 273 -200
rect 273 -201 274 -200
rect 274 -201 275 -200
rect 275 -201 276 -200
rect 276 -201 277 -200
rect 277 -201 278 -200
rect 278 -201 279 -200
rect 279 -201 280 -200
rect 280 -201 281 -200
rect 281 -201 282 -200
rect 282 -201 283 -200
rect 283 -201 284 -200
rect 284 -201 285 -200
rect 285 -201 286 -200
rect 286 -201 287 -200
rect 287 -201 288 -200
rect 288 -201 289 -200
rect 289 -201 290 -200
rect 290 -201 291 -200
rect 291 -201 292 -200
rect 292 -201 293 -200
rect 293 -201 294 -200
rect 294 -201 295 -200
rect 295 -201 296 -200
rect 296 -201 297 -200
rect 297 -201 298 -200
rect 298 -201 299 -200
rect 299 -201 300 -200
rect 300 -201 301 -200
rect 301 -201 302 -200
rect 302 -201 303 -200
rect 303 -201 304 -200
rect 304 -201 305 -200
rect 305 -201 306 -200
rect 306 -201 307 -200
rect 307 -201 308 -200
rect 308 -201 309 -200
rect 309 -201 310 -200
rect 310 -201 311 -200
rect 311 -201 312 -200
rect 312 -201 313 -200
rect 313 -201 314 -200
rect 314 -201 315 -200
rect 315 -201 316 -200
rect 316 -201 317 -200
rect 317 -201 318 -200
rect 318 -201 319 -200
rect 319 -201 320 -200
rect 320 -201 321 -200
rect 321 -201 322 -200
rect 322 -201 323 -200
rect 323 -201 324 -200
rect 324 -201 325 -200
rect 325 -201 326 -200
rect 326 -201 327 -200
rect 327 -201 328 -200
rect 328 -201 329 -200
rect 329 -201 330 -200
rect 330 -201 331 -200
rect 331 -201 332 -200
rect 332 -201 333 -200
rect 333 -201 334 -200
rect 334 -201 335 -200
rect 335 -201 336 -200
rect 336 -201 337 -200
rect 337 -201 338 -200
rect 338 -201 339 -200
rect 339 -201 340 -200
rect 340 -201 341 -200
rect 341 -201 342 -200
rect 342 -201 343 -200
rect 343 -201 344 -200
rect 344 -201 345 -200
rect 345 -201 346 -200
rect 346 -201 347 -200
rect 347 -201 348 -200
rect 348 -201 349 -200
rect 349 -201 350 -200
rect 350 -201 351 -200
rect 351 -201 352 -200
rect 352 -201 353 -200
rect 353 -201 354 -200
rect 354 -201 355 -200
rect 355 -201 356 -200
rect 356 -201 357 -200
rect 357 -201 358 -200
rect 358 -201 359 -200
rect 359 -201 360 -200
rect 360 -201 361 -200
rect 361 -201 362 -200
rect 362 -201 363 -200
rect 363 -201 364 -200
rect 364 -201 365 -200
rect 365 -201 366 -200
rect 366 -201 367 -200
rect 367 -201 368 -200
rect 368 -201 369 -200
rect 369 -201 370 -200
rect 370 -201 371 -200
rect 371 -201 372 -200
rect 372 -201 373 -200
rect 373 -201 374 -200
rect 374 -201 375 -200
rect 375 -201 376 -200
rect 376 -201 377 -200
rect 377 -201 378 -200
rect 378 -201 379 -200
rect 379 -201 380 -200
rect 380 -201 381 -200
rect 381 -201 382 -200
rect 382 -201 383 -200
rect 383 -201 384 -200
rect 384 -201 385 -200
rect 385 -201 386 -200
rect 386 -201 387 -200
rect 387 -201 388 -200
rect 388 -201 389 -200
rect 389 -201 390 -200
rect 390 -201 391 -200
rect 391 -201 392 -200
rect 392 -201 393 -200
rect 393 -201 394 -200
rect 394 -201 395 -200
rect 395 -201 396 -200
rect 396 -201 397 -200
rect 397 -201 398 -200
rect 398 -201 399 -200
rect 399 -201 400 -200
rect 400 -201 401 -200
rect 401 -201 402 -200
rect 402 -201 403 -200
rect 403 -201 404 -200
rect 404 -201 405 -200
rect 405 -201 406 -200
rect 406 -201 407 -200
rect 407 -201 408 -200
rect 408 -201 409 -200
rect 409 -201 410 -200
rect 410 -201 411 -200
rect 411 -201 412 -200
rect 412 -201 413 -200
rect 413 -201 414 -200
rect 414 -201 415 -200
rect 415 -201 416 -200
rect 416 -201 417 -200
rect 417 -201 418 -200
rect 418 -201 419 -200
rect 419 -201 420 -200
rect 420 -201 421 -200
rect 421 -201 422 -200
rect 422 -201 423 -200
rect 423 -201 424 -200
rect 424 -201 425 -200
rect 425 -201 426 -200
rect 426 -201 427 -200
rect 427 -201 428 -200
rect 428 -201 429 -200
rect 429 -201 430 -200
rect 430 -201 431 -200
rect 431 -201 432 -200
rect 432 -201 433 -200
rect 433 -201 434 -200
rect 434 -201 435 -200
rect 435 -201 436 -200
rect 436 -201 437 -200
rect 437 -201 438 -200
rect 438 -201 439 -200
rect 439 -201 440 -200
rect 440 -201 441 -200
rect 441 -201 442 -200
rect 442 -201 443 -200
rect 443 -201 444 -200
rect 444 -201 445 -200
rect 445 -201 446 -200
rect 446 -201 447 -200
rect 447 -201 448 -200
rect 448 -201 449 -200
rect 449 -201 450 -200
rect 450 -201 451 -200
rect 451 -201 452 -200
rect 452 -201 453 -200
rect 453 -201 454 -200
rect 454 -201 455 -200
rect 455 -201 456 -200
rect 456 -201 457 -200
rect 457 -201 458 -200
rect 458 -201 459 -200
rect 459 -201 460 -200
rect 460 -201 461 -200
rect 461 -201 462 -200
rect 462 -201 463 -200
rect 463 -201 464 -200
rect 464 -201 465 -200
rect 465 -201 466 -200
rect 466 -201 467 -200
rect 467 -201 468 -200
rect 468 -201 469 -200
rect 469 -201 470 -200
rect 470 -201 471 -200
rect 471 -201 472 -200
rect 472 -201 473 -200
rect 473 -201 474 -200
rect 474 -201 475 -200
rect 475 -201 476 -200
rect 476 -201 477 -200
rect 477 -201 478 -200
rect 478 -201 479 -200
rect 479 -201 480 -200
rect 2 -202 3 -201
rect 3 -202 4 -201
rect 4 -202 5 -201
rect 5 -202 6 -201
rect 6 -202 7 -201
rect 7 -202 8 -201
rect 8 -202 9 -201
rect 9 -202 10 -201
rect 10 -202 11 -201
rect 11 -202 12 -201
rect 12 -202 13 -201
rect 13 -202 14 -201
rect 14 -202 15 -201
rect 15 -202 16 -201
rect 16 -202 17 -201
rect 17 -202 18 -201
rect 18 -202 19 -201
rect 19 -202 20 -201
rect 20 -202 21 -201
rect 21 -202 22 -201
rect 22 -202 23 -201
rect 23 -202 24 -201
rect 24 -202 25 -201
rect 25 -202 26 -201
rect 26 -202 27 -201
rect 27 -202 28 -201
rect 28 -202 29 -201
rect 29 -202 30 -201
rect 30 -202 31 -201
rect 31 -202 32 -201
rect 32 -202 33 -201
rect 33 -202 34 -201
rect 34 -202 35 -201
rect 35 -202 36 -201
rect 36 -202 37 -201
rect 37 -202 38 -201
rect 38 -202 39 -201
rect 39 -202 40 -201
rect 40 -202 41 -201
rect 41 -202 42 -201
rect 42 -202 43 -201
rect 43 -202 44 -201
rect 44 -202 45 -201
rect 45 -202 46 -201
rect 46 -202 47 -201
rect 47 -202 48 -201
rect 48 -202 49 -201
rect 49 -202 50 -201
rect 50 -202 51 -201
rect 51 -202 52 -201
rect 52 -202 53 -201
rect 53 -202 54 -201
rect 54 -202 55 -201
rect 55 -202 56 -201
rect 56 -202 57 -201
rect 57 -202 58 -201
rect 58 -202 59 -201
rect 59 -202 60 -201
rect 60 -202 61 -201
rect 61 -202 62 -201
rect 62 -202 63 -201
rect 63 -202 64 -201
rect 64 -202 65 -201
rect 65 -202 66 -201
rect 66 -202 67 -201
rect 67 -202 68 -201
rect 68 -202 69 -201
rect 69 -202 70 -201
rect 70 -202 71 -201
rect 71 -202 72 -201
rect 72 -202 73 -201
rect 73 -202 74 -201
rect 74 -202 75 -201
rect 75 -202 76 -201
rect 76 -202 77 -201
rect 77 -202 78 -201
rect 78 -202 79 -201
rect 79 -202 80 -201
rect 80 -202 81 -201
rect 81 -202 82 -201
rect 82 -202 83 -201
rect 83 -202 84 -201
rect 84 -202 85 -201
rect 85 -202 86 -201
rect 86 -202 87 -201
rect 87 -202 88 -201
rect 88 -202 89 -201
rect 89 -202 90 -201
rect 90 -202 91 -201
rect 91 -202 92 -201
rect 92 -202 93 -201
rect 93 -202 94 -201
rect 94 -202 95 -201
rect 95 -202 96 -201
rect 96 -202 97 -201
rect 97 -202 98 -201
rect 98 -202 99 -201
rect 99 -202 100 -201
rect 100 -202 101 -201
rect 101 -202 102 -201
rect 102 -202 103 -201
rect 103 -202 104 -201
rect 104 -202 105 -201
rect 105 -202 106 -201
rect 106 -202 107 -201
rect 107 -202 108 -201
rect 108 -202 109 -201
rect 109 -202 110 -201
rect 110 -202 111 -201
rect 111 -202 112 -201
rect 112 -202 113 -201
rect 113 -202 114 -201
rect 114 -202 115 -201
rect 115 -202 116 -201
rect 116 -202 117 -201
rect 117 -202 118 -201
rect 118 -202 119 -201
rect 119 -202 120 -201
rect 120 -202 121 -201
rect 121 -202 122 -201
rect 122 -202 123 -201
rect 123 -202 124 -201
rect 124 -202 125 -201
rect 125 -202 126 -201
rect 126 -202 127 -201
rect 127 -202 128 -201
rect 128 -202 129 -201
rect 129 -202 130 -201
rect 130 -202 131 -201
rect 131 -202 132 -201
rect 132 -202 133 -201
rect 133 -202 134 -201
rect 134 -202 135 -201
rect 135 -202 136 -201
rect 136 -202 137 -201
rect 137 -202 138 -201
rect 138 -202 139 -201
rect 139 -202 140 -201
rect 140 -202 141 -201
rect 141 -202 142 -201
rect 142 -202 143 -201
rect 143 -202 144 -201
rect 144 -202 145 -201
rect 145 -202 146 -201
rect 146 -202 147 -201
rect 147 -202 148 -201
rect 148 -202 149 -201
rect 149 -202 150 -201
rect 150 -202 151 -201
rect 151 -202 152 -201
rect 152 -202 153 -201
rect 153 -202 154 -201
rect 154 -202 155 -201
rect 155 -202 156 -201
rect 156 -202 157 -201
rect 157 -202 158 -201
rect 158 -202 159 -201
rect 159 -202 160 -201
rect 160 -202 161 -201
rect 161 -202 162 -201
rect 162 -202 163 -201
rect 163 -202 164 -201
rect 164 -202 165 -201
rect 165 -202 166 -201
rect 166 -202 167 -201
rect 167 -202 168 -201
rect 168 -202 169 -201
rect 169 -202 170 -201
rect 170 -202 171 -201
rect 171 -202 172 -201
rect 172 -202 173 -201
rect 173 -202 174 -201
rect 174 -202 175 -201
rect 175 -202 176 -201
rect 176 -202 177 -201
rect 177 -202 178 -201
rect 178 -202 179 -201
rect 179 -202 180 -201
rect 180 -202 181 -201
rect 181 -202 182 -201
rect 182 -202 183 -201
rect 183 -202 184 -201
rect 184 -202 185 -201
rect 185 -202 186 -201
rect 186 -202 187 -201
rect 187 -202 188 -201
rect 188 -202 189 -201
rect 189 -202 190 -201
rect 190 -202 191 -201
rect 191 -202 192 -201
rect 192 -202 193 -201
rect 193 -202 194 -201
rect 194 -202 195 -201
rect 195 -202 196 -201
rect 196 -202 197 -201
rect 197 -202 198 -201
rect 198 -202 199 -201
rect 199 -202 200 -201
rect 200 -202 201 -201
rect 201 -202 202 -201
rect 202 -202 203 -201
rect 203 -202 204 -201
rect 204 -202 205 -201
rect 205 -202 206 -201
rect 206 -202 207 -201
rect 207 -202 208 -201
rect 208 -202 209 -201
rect 209 -202 210 -201
rect 210 -202 211 -201
rect 211 -202 212 -201
rect 212 -202 213 -201
rect 213 -202 214 -201
rect 214 -202 215 -201
rect 215 -202 216 -201
rect 216 -202 217 -201
rect 217 -202 218 -201
rect 218 -202 219 -201
rect 219 -202 220 -201
rect 220 -202 221 -201
rect 221 -202 222 -201
rect 222 -202 223 -201
rect 223 -202 224 -201
rect 224 -202 225 -201
rect 225 -202 226 -201
rect 226 -202 227 -201
rect 227 -202 228 -201
rect 228 -202 229 -201
rect 229 -202 230 -201
rect 230 -202 231 -201
rect 231 -202 232 -201
rect 232 -202 233 -201
rect 233 -202 234 -201
rect 234 -202 235 -201
rect 235 -202 236 -201
rect 236 -202 237 -201
rect 237 -202 238 -201
rect 238 -202 239 -201
rect 239 -202 240 -201
rect 240 -202 241 -201
rect 241 -202 242 -201
rect 242 -202 243 -201
rect 243 -202 244 -201
rect 244 -202 245 -201
rect 245 -202 246 -201
rect 246 -202 247 -201
rect 247 -202 248 -201
rect 248 -202 249 -201
rect 249 -202 250 -201
rect 250 -202 251 -201
rect 251 -202 252 -201
rect 252 -202 253 -201
rect 253 -202 254 -201
rect 254 -202 255 -201
rect 255 -202 256 -201
rect 256 -202 257 -201
rect 257 -202 258 -201
rect 258 -202 259 -201
rect 259 -202 260 -201
rect 260 -202 261 -201
rect 261 -202 262 -201
rect 262 -202 263 -201
rect 263 -202 264 -201
rect 264 -202 265 -201
rect 265 -202 266 -201
rect 266 -202 267 -201
rect 267 -202 268 -201
rect 268 -202 269 -201
rect 269 -202 270 -201
rect 270 -202 271 -201
rect 271 -202 272 -201
rect 272 -202 273 -201
rect 273 -202 274 -201
rect 274 -202 275 -201
rect 275 -202 276 -201
rect 276 -202 277 -201
rect 277 -202 278 -201
rect 278 -202 279 -201
rect 279 -202 280 -201
rect 280 -202 281 -201
rect 281 -202 282 -201
rect 282 -202 283 -201
rect 283 -202 284 -201
rect 284 -202 285 -201
rect 285 -202 286 -201
rect 286 -202 287 -201
rect 287 -202 288 -201
rect 288 -202 289 -201
rect 289 -202 290 -201
rect 290 -202 291 -201
rect 291 -202 292 -201
rect 292 -202 293 -201
rect 293 -202 294 -201
rect 294 -202 295 -201
rect 295 -202 296 -201
rect 296 -202 297 -201
rect 297 -202 298 -201
rect 298 -202 299 -201
rect 299 -202 300 -201
rect 300 -202 301 -201
rect 301 -202 302 -201
rect 302 -202 303 -201
rect 303 -202 304 -201
rect 304 -202 305 -201
rect 305 -202 306 -201
rect 306 -202 307 -201
rect 307 -202 308 -201
rect 308 -202 309 -201
rect 309 -202 310 -201
rect 310 -202 311 -201
rect 311 -202 312 -201
rect 312 -202 313 -201
rect 313 -202 314 -201
rect 314 -202 315 -201
rect 315 -202 316 -201
rect 316 -202 317 -201
rect 317 -202 318 -201
rect 318 -202 319 -201
rect 319 -202 320 -201
rect 320 -202 321 -201
rect 321 -202 322 -201
rect 322 -202 323 -201
rect 323 -202 324 -201
rect 324 -202 325 -201
rect 325 -202 326 -201
rect 326 -202 327 -201
rect 327 -202 328 -201
rect 328 -202 329 -201
rect 329 -202 330 -201
rect 330 -202 331 -201
rect 331 -202 332 -201
rect 332 -202 333 -201
rect 333 -202 334 -201
rect 334 -202 335 -201
rect 335 -202 336 -201
rect 336 -202 337 -201
rect 337 -202 338 -201
rect 338 -202 339 -201
rect 339 -202 340 -201
rect 340 -202 341 -201
rect 341 -202 342 -201
rect 342 -202 343 -201
rect 343 -202 344 -201
rect 344 -202 345 -201
rect 345 -202 346 -201
rect 346 -202 347 -201
rect 347 -202 348 -201
rect 348 -202 349 -201
rect 349 -202 350 -201
rect 350 -202 351 -201
rect 351 -202 352 -201
rect 352 -202 353 -201
rect 353 -202 354 -201
rect 354 -202 355 -201
rect 355 -202 356 -201
rect 356 -202 357 -201
rect 357 -202 358 -201
rect 358 -202 359 -201
rect 359 -202 360 -201
rect 360 -202 361 -201
rect 361 -202 362 -201
rect 362 -202 363 -201
rect 363 -202 364 -201
rect 364 -202 365 -201
rect 365 -202 366 -201
rect 366 -202 367 -201
rect 367 -202 368 -201
rect 368 -202 369 -201
rect 369 -202 370 -201
rect 370 -202 371 -201
rect 371 -202 372 -201
rect 372 -202 373 -201
rect 373 -202 374 -201
rect 374 -202 375 -201
rect 375 -202 376 -201
rect 376 -202 377 -201
rect 377 -202 378 -201
rect 378 -202 379 -201
rect 379 -202 380 -201
rect 380 -202 381 -201
rect 381 -202 382 -201
rect 382 -202 383 -201
rect 383 -202 384 -201
rect 384 -202 385 -201
rect 385 -202 386 -201
rect 386 -202 387 -201
rect 387 -202 388 -201
rect 388 -202 389 -201
rect 389 -202 390 -201
rect 390 -202 391 -201
rect 391 -202 392 -201
rect 392 -202 393 -201
rect 393 -202 394 -201
rect 394 -202 395 -201
rect 395 -202 396 -201
rect 396 -202 397 -201
rect 397 -202 398 -201
rect 398 -202 399 -201
rect 399 -202 400 -201
rect 400 -202 401 -201
rect 401 -202 402 -201
rect 402 -202 403 -201
rect 403 -202 404 -201
rect 404 -202 405 -201
rect 405 -202 406 -201
rect 406 -202 407 -201
rect 407 -202 408 -201
rect 408 -202 409 -201
rect 409 -202 410 -201
rect 410 -202 411 -201
rect 411 -202 412 -201
rect 412 -202 413 -201
rect 413 -202 414 -201
rect 414 -202 415 -201
rect 415 -202 416 -201
rect 416 -202 417 -201
rect 417 -202 418 -201
rect 418 -202 419 -201
rect 419 -202 420 -201
rect 420 -202 421 -201
rect 421 -202 422 -201
rect 422 -202 423 -201
rect 423 -202 424 -201
rect 424 -202 425 -201
rect 425 -202 426 -201
rect 426 -202 427 -201
rect 427 -202 428 -201
rect 428 -202 429 -201
rect 429 -202 430 -201
rect 430 -202 431 -201
rect 431 -202 432 -201
rect 432 -202 433 -201
rect 433 -202 434 -201
rect 434 -202 435 -201
rect 435 -202 436 -201
rect 436 -202 437 -201
rect 437 -202 438 -201
rect 438 -202 439 -201
rect 439 -202 440 -201
rect 440 -202 441 -201
rect 441 -202 442 -201
rect 442 -202 443 -201
rect 443 -202 444 -201
rect 444 -202 445 -201
rect 445 -202 446 -201
rect 446 -202 447 -201
rect 447 -202 448 -201
rect 448 -202 449 -201
rect 449 -202 450 -201
rect 450 -202 451 -201
rect 451 -202 452 -201
rect 452 -202 453 -201
rect 453 -202 454 -201
rect 454 -202 455 -201
rect 455 -202 456 -201
rect 456 -202 457 -201
rect 457 -202 458 -201
rect 458 -202 459 -201
rect 459 -202 460 -201
rect 460 -202 461 -201
rect 461 -202 462 -201
rect 462 -202 463 -201
rect 463 -202 464 -201
rect 464 -202 465 -201
rect 465 -202 466 -201
rect 466 -202 467 -201
rect 467 -202 468 -201
rect 468 -202 469 -201
rect 469 -202 470 -201
rect 470 -202 471 -201
rect 471 -202 472 -201
rect 472 -202 473 -201
rect 473 -202 474 -201
rect 474 -202 475 -201
rect 475 -202 476 -201
rect 476 -202 477 -201
rect 477 -202 478 -201
rect 478 -202 479 -201
rect 479 -202 480 -201
rect 2 -203 3 -202
rect 3 -203 4 -202
rect 4 -203 5 -202
rect 5 -203 6 -202
rect 6 -203 7 -202
rect 7 -203 8 -202
rect 8 -203 9 -202
rect 9 -203 10 -202
rect 10 -203 11 -202
rect 11 -203 12 -202
rect 12 -203 13 -202
rect 13 -203 14 -202
rect 14 -203 15 -202
rect 15 -203 16 -202
rect 16 -203 17 -202
rect 17 -203 18 -202
rect 18 -203 19 -202
rect 19 -203 20 -202
rect 20 -203 21 -202
rect 21 -203 22 -202
rect 22 -203 23 -202
rect 23 -203 24 -202
rect 24 -203 25 -202
rect 25 -203 26 -202
rect 26 -203 27 -202
rect 27 -203 28 -202
rect 28 -203 29 -202
rect 29 -203 30 -202
rect 30 -203 31 -202
rect 31 -203 32 -202
rect 32 -203 33 -202
rect 33 -203 34 -202
rect 34 -203 35 -202
rect 35 -203 36 -202
rect 36 -203 37 -202
rect 37 -203 38 -202
rect 38 -203 39 -202
rect 39 -203 40 -202
rect 40 -203 41 -202
rect 41 -203 42 -202
rect 42 -203 43 -202
rect 43 -203 44 -202
rect 44 -203 45 -202
rect 45 -203 46 -202
rect 46 -203 47 -202
rect 47 -203 48 -202
rect 48 -203 49 -202
rect 49 -203 50 -202
rect 50 -203 51 -202
rect 51 -203 52 -202
rect 52 -203 53 -202
rect 53 -203 54 -202
rect 54 -203 55 -202
rect 55 -203 56 -202
rect 56 -203 57 -202
rect 57 -203 58 -202
rect 58 -203 59 -202
rect 59 -203 60 -202
rect 60 -203 61 -202
rect 61 -203 62 -202
rect 62 -203 63 -202
rect 63 -203 64 -202
rect 64 -203 65 -202
rect 65 -203 66 -202
rect 66 -203 67 -202
rect 67 -203 68 -202
rect 68 -203 69 -202
rect 69 -203 70 -202
rect 70 -203 71 -202
rect 71 -203 72 -202
rect 72 -203 73 -202
rect 73 -203 74 -202
rect 74 -203 75 -202
rect 75 -203 76 -202
rect 76 -203 77 -202
rect 77 -203 78 -202
rect 78 -203 79 -202
rect 79 -203 80 -202
rect 80 -203 81 -202
rect 81 -203 82 -202
rect 82 -203 83 -202
rect 83 -203 84 -202
rect 84 -203 85 -202
rect 85 -203 86 -202
rect 86 -203 87 -202
rect 87 -203 88 -202
rect 88 -203 89 -202
rect 89 -203 90 -202
rect 90 -203 91 -202
rect 91 -203 92 -202
rect 92 -203 93 -202
rect 93 -203 94 -202
rect 94 -203 95 -202
rect 95 -203 96 -202
rect 96 -203 97 -202
rect 97 -203 98 -202
rect 98 -203 99 -202
rect 99 -203 100 -202
rect 100 -203 101 -202
rect 101 -203 102 -202
rect 102 -203 103 -202
rect 103 -203 104 -202
rect 104 -203 105 -202
rect 105 -203 106 -202
rect 106 -203 107 -202
rect 107 -203 108 -202
rect 108 -203 109 -202
rect 109 -203 110 -202
rect 110 -203 111 -202
rect 111 -203 112 -202
rect 112 -203 113 -202
rect 113 -203 114 -202
rect 114 -203 115 -202
rect 115 -203 116 -202
rect 116 -203 117 -202
rect 117 -203 118 -202
rect 118 -203 119 -202
rect 119 -203 120 -202
rect 120 -203 121 -202
rect 121 -203 122 -202
rect 122 -203 123 -202
rect 123 -203 124 -202
rect 124 -203 125 -202
rect 125 -203 126 -202
rect 126 -203 127 -202
rect 127 -203 128 -202
rect 128 -203 129 -202
rect 129 -203 130 -202
rect 130 -203 131 -202
rect 131 -203 132 -202
rect 132 -203 133 -202
rect 133 -203 134 -202
rect 134 -203 135 -202
rect 135 -203 136 -202
rect 136 -203 137 -202
rect 137 -203 138 -202
rect 138 -203 139 -202
rect 139 -203 140 -202
rect 140 -203 141 -202
rect 141 -203 142 -202
rect 142 -203 143 -202
rect 143 -203 144 -202
rect 144 -203 145 -202
rect 145 -203 146 -202
rect 146 -203 147 -202
rect 147 -203 148 -202
rect 148 -203 149 -202
rect 149 -203 150 -202
rect 150 -203 151 -202
rect 151 -203 152 -202
rect 152 -203 153 -202
rect 153 -203 154 -202
rect 154 -203 155 -202
rect 155 -203 156 -202
rect 156 -203 157 -202
rect 157 -203 158 -202
rect 158 -203 159 -202
rect 159 -203 160 -202
rect 160 -203 161 -202
rect 161 -203 162 -202
rect 162 -203 163 -202
rect 163 -203 164 -202
rect 164 -203 165 -202
rect 165 -203 166 -202
rect 166 -203 167 -202
rect 167 -203 168 -202
rect 168 -203 169 -202
rect 169 -203 170 -202
rect 170 -203 171 -202
rect 171 -203 172 -202
rect 172 -203 173 -202
rect 173 -203 174 -202
rect 174 -203 175 -202
rect 175 -203 176 -202
rect 176 -203 177 -202
rect 177 -203 178 -202
rect 178 -203 179 -202
rect 179 -203 180 -202
rect 180 -203 181 -202
rect 181 -203 182 -202
rect 182 -203 183 -202
rect 183 -203 184 -202
rect 184 -203 185 -202
rect 185 -203 186 -202
rect 186 -203 187 -202
rect 187 -203 188 -202
rect 188 -203 189 -202
rect 189 -203 190 -202
rect 190 -203 191 -202
rect 191 -203 192 -202
rect 192 -203 193 -202
rect 193 -203 194 -202
rect 194 -203 195 -202
rect 195 -203 196 -202
rect 196 -203 197 -202
rect 197 -203 198 -202
rect 198 -203 199 -202
rect 199 -203 200 -202
rect 200 -203 201 -202
rect 201 -203 202 -202
rect 202 -203 203 -202
rect 203 -203 204 -202
rect 204 -203 205 -202
rect 205 -203 206 -202
rect 206 -203 207 -202
rect 207 -203 208 -202
rect 208 -203 209 -202
rect 209 -203 210 -202
rect 210 -203 211 -202
rect 211 -203 212 -202
rect 212 -203 213 -202
rect 213 -203 214 -202
rect 214 -203 215 -202
rect 215 -203 216 -202
rect 216 -203 217 -202
rect 217 -203 218 -202
rect 218 -203 219 -202
rect 219 -203 220 -202
rect 220 -203 221 -202
rect 221 -203 222 -202
rect 222 -203 223 -202
rect 223 -203 224 -202
rect 224 -203 225 -202
rect 225 -203 226 -202
rect 226 -203 227 -202
rect 227 -203 228 -202
rect 228 -203 229 -202
rect 229 -203 230 -202
rect 230 -203 231 -202
rect 231 -203 232 -202
rect 232 -203 233 -202
rect 233 -203 234 -202
rect 234 -203 235 -202
rect 235 -203 236 -202
rect 236 -203 237 -202
rect 237 -203 238 -202
rect 238 -203 239 -202
rect 239 -203 240 -202
rect 240 -203 241 -202
rect 241 -203 242 -202
rect 242 -203 243 -202
rect 243 -203 244 -202
rect 244 -203 245 -202
rect 245 -203 246 -202
rect 246 -203 247 -202
rect 247 -203 248 -202
rect 248 -203 249 -202
rect 249 -203 250 -202
rect 250 -203 251 -202
rect 251 -203 252 -202
rect 252 -203 253 -202
rect 253 -203 254 -202
rect 254 -203 255 -202
rect 255 -203 256 -202
rect 256 -203 257 -202
rect 257 -203 258 -202
rect 258 -203 259 -202
rect 259 -203 260 -202
rect 260 -203 261 -202
rect 261 -203 262 -202
rect 262 -203 263 -202
rect 263 -203 264 -202
rect 264 -203 265 -202
rect 265 -203 266 -202
rect 266 -203 267 -202
rect 267 -203 268 -202
rect 268 -203 269 -202
rect 269 -203 270 -202
rect 270 -203 271 -202
rect 271 -203 272 -202
rect 272 -203 273 -202
rect 273 -203 274 -202
rect 274 -203 275 -202
rect 275 -203 276 -202
rect 276 -203 277 -202
rect 277 -203 278 -202
rect 278 -203 279 -202
rect 279 -203 280 -202
rect 280 -203 281 -202
rect 281 -203 282 -202
rect 282 -203 283 -202
rect 283 -203 284 -202
rect 284 -203 285 -202
rect 285 -203 286 -202
rect 286 -203 287 -202
rect 287 -203 288 -202
rect 288 -203 289 -202
rect 289 -203 290 -202
rect 290 -203 291 -202
rect 291 -203 292 -202
rect 292 -203 293 -202
rect 293 -203 294 -202
rect 294 -203 295 -202
rect 295 -203 296 -202
rect 296 -203 297 -202
rect 297 -203 298 -202
rect 298 -203 299 -202
rect 299 -203 300 -202
rect 300 -203 301 -202
rect 301 -203 302 -202
rect 302 -203 303 -202
rect 303 -203 304 -202
rect 304 -203 305 -202
rect 305 -203 306 -202
rect 306 -203 307 -202
rect 307 -203 308 -202
rect 308 -203 309 -202
rect 309 -203 310 -202
rect 310 -203 311 -202
rect 311 -203 312 -202
rect 312 -203 313 -202
rect 313 -203 314 -202
rect 314 -203 315 -202
rect 315 -203 316 -202
rect 316 -203 317 -202
rect 317 -203 318 -202
rect 318 -203 319 -202
rect 319 -203 320 -202
rect 320 -203 321 -202
rect 321 -203 322 -202
rect 322 -203 323 -202
rect 323 -203 324 -202
rect 324 -203 325 -202
rect 325 -203 326 -202
rect 326 -203 327 -202
rect 327 -203 328 -202
rect 328 -203 329 -202
rect 329 -203 330 -202
rect 330 -203 331 -202
rect 331 -203 332 -202
rect 332 -203 333 -202
rect 333 -203 334 -202
rect 334 -203 335 -202
rect 335 -203 336 -202
rect 336 -203 337 -202
rect 337 -203 338 -202
rect 338 -203 339 -202
rect 339 -203 340 -202
rect 340 -203 341 -202
rect 341 -203 342 -202
rect 342 -203 343 -202
rect 343 -203 344 -202
rect 344 -203 345 -202
rect 345 -203 346 -202
rect 346 -203 347 -202
rect 347 -203 348 -202
rect 348 -203 349 -202
rect 349 -203 350 -202
rect 350 -203 351 -202
rect 351 -203 352 -202
rect 352 -203 353 -202
rect 353 -203 354 -202
rect 354 -203 355 -202
rect 355 -203 356 -202
rect 356 -203 357 -202
rect 357 -203 358 -202
rect 358 -203 359 -202
rect 359 -203 360 -202
rect 360 -203 361 -202
rect 361 -203 362 -202
rect 362 -203 363 -202
rect 363 -203 364 -202
rect 364 -203 365 -202
rect 365 -203 366 -202
rect 366 -203 367 -202
rect 367 -203 368 -202
rect 368 -203 369 -202
rect 369 -203 370 -202
rect 370 -203 371 -202
rect 371 -203 372 -202
rect 372 -203 373 -202
rect 373 -203 374 -202
rect 374 -203 375 -202
rect 375 -203 376 -202
rect 376 -203 377 -202
rect 377 -203 378 -202
rect 378 -203 379 -202
rect 379 -203 380 -202
rect 380 -203 381 -202
rect 381 -203 382 -202
rect 382 -203 383 -202
rect 383 -203 384 -202
rect 384 -203 385 -202
rect 385 -203 386 -202
rect 386 -203 387 -202
rect 387 -203 388 -202
rect 388 -203 389 -202
rect 389 -203 390 -202
rect 390 -203 391 -202
rect 391 -203 392 -202
rect 392 -203 393 -202
rect 393 -203 394 -202
rect 394 -203 395 -202
rect 395 -203 396 -202
rect 396 -203 397 -202
rect 397 -203 398 -202
rect 398 -203 399 -202
rect 399 -203 400 -202
rect 400 -203 401 -202
rect 401 -203 402 -202
rect 402 -203 403 -202
rect 403 -203 404 -202
rect 404 -203 405 -202
rect 405 -203 406 -202
rect 406 -203 407 -202
rect 407 -203 408 -202
rect 408 -203 409 -202
rect 409 -203 410 -202
rect 410 -203 411 -202
rect 411 -203 412 -202
rect 412 -203 413 -202
rect 413 -203 414 -202
rect 414 -203 415 -202
rect 415 -203 416 -202
rect 416 -203 417 -202
rect 417 -203 418 -202
rect 418 -203 419 -202
rect 419 -203 420 -202
rect 420 -203 421 -202
rect 421 -203 422 -202
rect 422 -203 423 -202
rect 423 -203 424 -202
rect 424 -203 425 -202
rect 425 -203 426 -202
rect 426 -203 427 -202
rect 427 -203 428 -202
rect 428 -203 429 -202
rect 429 -203 430 -202
rect 430 -203 431 -202
rect 431 -203 432 -202
rect 432 -203 433 -202
rect 433 -203 434 -202
rect 434 -203 435 -202
rect 435 -203 436 -202
rect 436 -203 437 -202
rect 437 -203 438 -202
rect 438 -203 439 -202
rect 439 -203 440 -202
rect 440 -203 441 -202
rect 441 -203 442 -202
rect 442 -203 443 -202
rect 443 -203 444 -202
rect 444 -203 445 -202
rect 445 -203 446 -202
rect 446 -203 447 -202
rect 447 -203 448 -202
rect 448 -203 449 -202
rect 449 -203 450 -202
rect 450 -203 451 -202
rect 451 -203 452 -202
rect 452 -203 453 -202
rect 453 -203 454 -202
rect 454 -203 455 -202
rect 455 -203 456 -202
rect 456 -203 457 -202
rect 457 -203 458 -202
rect 458 -203 459 -202
rect 459 -203 460 -202
rect 460 -203 461 -202
rect 461 -203 462 -202
rect 462 -203 463 -202
rect 463 -203 464 -202
rect 464 -203 465 -202
rect 465 -203 466 -202
rect 466 -203 467 -202
rect 467 -203 468 -202
rect 468 -203 469 -202
rect 469 -203 470 -202
rect 470 -203 471 -202
rect 471 -203 472 -202
rect 472 -203 473 -202
rect 473 -203 474 -202
rect 474 -203 475 -202
rect 475 -203 476 -202
rect 476 -203 477 -202
rect 477 -203 478 -202
rect 478 -203 479 -202
rect 479 -203 480 -202
rect 2 -204 3 -203
rect 3 -204 4 -203
rect 4 -204 5 -203
rect 5 -204 6 -203
rect 6 -204 7 -203
rect 7 -204 8 -203
rect 8 -204 9 -203
rect 9 -204 10 -203
rect 10 -204 11 -203
rect 11 -204 12 -203
rect 12 -204 13 -203
rect 13 -204 14 -203
rect 14 -204 15 -203
rect 15 -204 16 -203
rect 16 -204 17 -203
rect 17 -204 18 -203
rect 18 -204 19 -203
rect 19 -204 20 -203
rect 20 -204 21 -203
rect 21 -204 22 -203
rect 22 -204 23 -203
rect 23 -204 24 -203
rect 24 -204 25 -203
rect 25 -204 26 -203
rect 26 -204 27 -203
rect 27 -204 28 -203
rect 28 -204 29 -203
rect 29 -204 30 -203
rect 30 -204 31 -203
rect 31 -204 32 -203
rect 32 -204 33 -203
rect 33 -204 34 -203
rect 34 -204 35 -203
rect 35 -204 36 -203
rect 36 -204 37 -203
rect 37 -204 38 -203
rect 38 -204 39 -203
rect 39 -204 40 -203
rect 40 -204 41 -203
rect 41 -204 42 -203
rect 42 -204 43 -203
rect 43 -204 44 -203
rect 44 -204 45 -203
rect 45 -204 46 -203
rect 46 -204 47 -203
rect 47 -204 48 -203
rect 48 -204 49 -203
rect 49 -204 50 -203
rect 50 -204 51 -203
rect 51 -204 52 -203
rect 52 -204 53 -203
rect 53 -204 54 -203
rect 54 -204 55 -203
rect 55 -204 56 -203
rect 56 -204 57 -203
rect 57 -204 58 -203
rect 58 -204 59 -203
rect 59 -204 60 -203
rect 60 -204 61 -203
rect 61 -204 62 -203
rect 62 -204 63 -203
rect 63 -204 64 -203
rect 64 -204 65 -203
rect 65 -204 66 -203
rect 66 -204 67 -203
rect 67 -204 68 -203
rect 68 -204 69 -203
rect 69 -204 70 -203
rect 70 -204 71 -203
rect 71 -204 72 -203
rect 72 -204 73 -203
rect 73 -204 74 -203
rect 74 -204 75 -203
rect 75 -204 76 -203
rect 76 -204 77 -203
rect 77 -204 78 -203
rect 78 -204 79 -203
rect 79 -204 80 -203
rect 80 -204 81 -203
rect 81 -204 82 -203
rect 82 -204 83 -203
rect 83 -204 84 -203
rect 84 -204 85 -203
rect 85 -204 86 -203
rect 86 -204 87 -203
rect 87 -204 88 -203
rect 88 -204 89 -203
rect 89 -204 90 -203
rect 90 -204 91 -203
rect 91 -204 92 -203
rect 92 -204 93 -203
rect 93 -204 94 -203
rect 94 -204 95 -203
rect 95 -204 96 -203
rect 96 -204 97 -203
rect 97 -204 98 -203
rect 98 -204 99 -203
rect 99 -204 100 -203
rect 100 -204 101 -203
rect 101 -204 102 -203
rect 102 -204 103 -203
rect 103 -204 104 -203
rect 104 -204 105 -203
rect 105 -204 106 -203
rect 106 -204 107 -203
rect 107 -204 108 -203
rect 108 -204 109 -203
rect 109 -204 110 -203
rect 110 -204 111 -203
rect 111 -204 112 -203
rect 112 -204 113 -203
rect 113 -204 114 -203
rect 114 -204 115 -203
rect 115 -204 116 -203
rect 116 -204 117 -203
rect 117 -204 118 -203
rect 118 -204 119 -203
rect 119 -204 120 -203
rect 120 -204 121 -203
rect 121 -204 122 -203
rect 122 -204 123 -203
rect 123 -204 124 -203
rect 124 -204 125 -203
rect 125 -204 126 -203
rect 126 -204 127 -203
rect 127 -204 128 -203
rect 128 -204 129 -203
rect 129 -204 130 -203
rect 130 -204 131 -203
rect 131 -204 132 -203
rect 132 -204 133 -203
rect 133 -204 134 -203
rect 134 -204 135 -203
rect 135 -204 136 -203
rect 136 -204 137 -203
rect 137 -204 138 -203
rect 138 -204 139 -203
rect 139 -204 140 -203
rect 140 -204 141 -203
rect 141 -204 142 -203
rect 142 -204 143 -203
rect 143 -204 144 -203
rect 144 -204 145 -203
rect 145 -204 146 -203
rect 146 -204 147 -203
rect 147 -204 148 -203
rect 148 -204 149 -203
rect 149 -204 150 -203
rect 150 -204 151 -203
rect 151 -204 152 -203
rect 152 -204 153 -203
rect 153 -204 154 -203
rect 154 -204 155 -203
rect 155 -204 156 -203
rect 156 -204 157 -203
rect 157 -204 158 -203
rect 158 -204 159 -203
rect 159 -204 160 -203
rect 160 -204 161 -203
rect 161 -204 162 -203
rect 162 -204 163 -203
rect 163 -204 164 -203
rect 164 -204 165 -203
rect 165 -204 166 -203
rect 166 -204 167 -203
rect 167 -204 168 -203
rect 168 -204 169 -203
rect 169 -204 170 -203
rect 170 -204 171 -203
rect 171 -204 172 -203
rect 172 -204 173 -203
rect 173 -204 174 -203
rect 174 -204 175 -203
rect 175 -204 176 -203
rect 176 -204 177 -203
rect 177 -204 178 -203
rect 178 -204 179 -203
rect 179 -204 180 -203
rect 180 -204 181 -203
rect 181 -204 182 -203
rect 182 -204 183 -203
rect 183 -204 184 -203
rect 184 -204 185 -203
rect 185 -204 186 -203
rect 186 -204 187 -203
rect 187 -204 188 -203
rect 188 -204 189 -203
rect 189 -204 190 -203
rect 190 -204 191 -203
rect 191 -204 192 -203
rect 192 -204 193 -203
rect 193 -204 194 -203
rect 194 -204 195 -203
rect 195 -204 196 -203
rect 196 -204 197 -203
rect 197 -204 198 -203
rect 198 -204 199 -203
rect 199 -204 200 -203
rect 200 -204 201 -203
rect 201 -204 202 -203
rect 202 -204 203 -203
rect 203 -204 204 -203
rect 204 -204 205 -203
rect 205 -204 206 -203
rect 206 -204 207 -203
rect 207 -204 208 -203
rect 208 -204 209 -203
rect 209 -204 210 -203
rect 210 -204 211 -203
rect 211 -204 212 -203
rect 212 -204 213 -203
rect 213 -204 214 -203
rect 214 -204 215 -203
rect 215 -204 216 -203
rect 216 -204 217 -203
rect 217 -204 218 -203
rect 218 -204 219 -203
rect 219 -204 220 -203
rect 220 -204 221 -203
rect 221 -204 222 -203
rect 222 -204 223 -203
rect 223 -204 224 -203
rect 224 -204 225 -203
rect 225 -204 226 -203
rect 226 -204 227 -203
rect 227 -204 228 -203
rect 228 -204 229 -203
rect 229 -204 230 -203
rect 230 -204 231 -203
rect 231 -204 232 -203
rect 232 -204 233 -203
rect 233 -204 234 -203
rect 234 -204 235 -203
rect 235 -204 236 -203
rect 236 -204 237 -203
rect 237 -204 238 -203
rect 238 -204 239 -203
rect 239 -204 240 -203
rect 240 -204 241 -203
rect 241 -204 242 -203
rect 242 -204 243 -203
rect 243 -204 244 -203
rect 244 -204 245 -203
rect 245 -204 246 -203
rect 246 -204 247 -203
rect 247 -204 248 -203
rect 248 -204 249 -203
rect 249 -204 250 -203
rect 250 -204 251 -203
rect 251 -204 252 -203
rect 252 -204 253 -203
rect 253 -204 254 -203
rect 254 -204 255 -203
rect 255 -204 256 -203
rect 256 -204 257 -203
rect 257 -204 258 -203
rect 258 -204 259 -203
rect 259 -204 260 -203
rect 260 -204 261 -203
rect 261 -204 262 -203
rect 262 -204 263 -203
rect 263 -204 264 -203
rect 264 -204 265 -203
rect 265 -204 266 -203
rect 266 -204 267 -203
rect 267 -204 268 -203
rect 268 -204 269 -203
rect 269 -204 270 -203
rect 270 -204 271 -203
rect 271 -204 272 -203
rect 272 -204 273 -203
rect 273 -204 274 -203
rect 274 -204 275 -203
rect 275 -204 276 -203
rect 276 -204 277 -203
rect 277 -204 278 -203
rect 278 -204 279 -203
rect 279 -204 280 -203
rect 280 -204 281 -203
rect 281 -204 282 -203
rect 282 -204 283 -203
rect 283 -204 284 -203
rect 284 -204 285 -203
rect 285 -204 286 -203
rect 286 -204 287 -203
rect 287 -204 288 -203
rect 288 -204 289 -203
rect 289 -204 290 -203
rect 290 -204 291 -203
rect 291 -204 292 -203
rect 292 -204 293 -203
rect 293 -204 294 -203
rect 294 -204 295 -203
rect 295 -204 296 -203
rect 296 -204 297 -203
rect 297 -204 298 -203
rect 298 -204 299 -203
rect 299 -204 300 -203
rect 300 -204 301 -203
rect 301 -204 302 -203
rect 302 -204 303 -203
rect 303 -204 304 -203
rect 304 -204 305 -203
rect 305 -204 306 -203
rect 306 -204 307 -203
rect 307 -204 308 -203
rect 308 -204 309 -203
rect 309 -204 310 -203
rect 310 -204 311 -203
rect 311 -204 312 -203
rect 312 -204 313 -203
rect 313 -204 314 -203
rect 314 -204 315 -203
rect 315 -204 316 -203
rect 316 -204 317 -203
rect 317 -204 318 -203
rect 318 -204 319 -203
rect 319 -204 320 -203
rect 320 -204 321 -203
rect 321 -204 322 -203
rect 322 -204 323 -203
rect 323 -204 324 -203
rect 324 -204 325 -203
rect 325 -204 326 -203
rect 326 -204 327 -203
rect 327 -204 328 -203
rect 328 -204 329 -203
rect 329 -204 330 -203
rect 330 -204 331 -203
rect 331 -204 332 -203
rect 332 -204 333 -203
rect 333 -204 334 -203
rect 334 -204 335 -203
rect 335 -204 336 -203
rect 336 -204 337 -203
rect 337 -204 338 -203
rect 338 -204 339 -203
rect 339 -204 340 -203
rect 340 -204 341 -203
rect 341 -204 342 -203
rect 342 -204 343 -203
rect 343 -204 344 -203
rect 344 -204 345 -203
rect 345 -204 346 -203
rect 346 -204 347 -203
rect 347 -204 348 -203
rect 348 -204 349 -203
rect 349 -204 350 -203
rect 350 -204 351 -203
rect 351 -204 352 -203
rect 352 -204 353 -203
rect 353 -204 354 -203
rect 354 -204 355 -203
rect 355 -204 356 -203
rect 356 -204 357 -203
rect 357 -204 358 -203
rect 358 -204 359 -203
rect 359 -204 360 -203
rect 360 -204 361 -203
rect 361 -204 362 -203
rect 362 -204 363 -203
rect 363 -204 364 -203
rect 364 -204 365 -203
rect 365 -204 366 -203
rect 366 -204 367 -203
rect 367 -204 368 -203
rect 368 -204 369 -203
rect 369 -204 370 -203
rect 370 -204 371 -203
rect 371 -204 372 -203
rect 372 -204 373 -203
rect 373 -204 374 -203
rect 374 -204 375 -203
rect 375 -204 376 -203
rect 376 -204 377 -203
rect 377 -204 378 -203
rect 378 -204 379 -203
rect 379 -204 380 -203
rect 380 -204 381 -203
rect 381 -204 382 -203
rect 382 -204 383 -203
rect 383 -204 384 -203
rect 384 -204 385 -203
rect 385 -204 386 -203
rect 386 -204 387 -203
rect 387 -204 388 -203
rect 388 -204 389 -203
rect 389 -204 390 -203
rect 390 -204 391 -203
rect 391 -204 392 -203
rect 392 -204 393 -203
rect 393 -204 394 -203
rect 394 -204 395 -203
rect 395 -204 396 -203
rect 396 -204 397 -203
rect 397 -204 398 -203
rect 398 -204 399 -203
rect 399 -204 400 -203
rect 400 -204 401 -203
rect 401 -204 402 -203
rect 402 -204 403 -203
rect 403 -204 404 -203
rect 404 -204 405 -203
rect 405 -204 406 -203
rect 406 -204 407 -203
rect 407 -204 408 -203
rect 408 -204 409 -203
rect 409 -204 410 -203
rect 410 -204 411 -203
rect 411 -204 412 -203
rect 412 -204 413 -203
rect 413 -204 414 -203
rect 414 -204 415 -203
rect 415 -204 416 -203
rect 416 -204 417 -203
rect 417 -204 418 -203
rect 418 -204 419 -203
rect 419 -204 420 -203
rect 420 -204 421 -203
rect 421 -204 422 -203
rect 422 -204 423 -203
rect 423 -204 424 -203
rect 424 -204 425 -203
rect 425 -204 426 -203
rect 426 -204 427 -203
rect 427 -204 428 -203
rect 428 -204 429 -203
rect 429 -204 430 -203
rect 430 -204 431 -203
rect 431 -204 432 -203
rect 432 -204 433 -203
rect 433 -204 434 -203
rect 434 -204 435 -203
rect 435 -204 436 -203
rect 436 -204 437 -203
rect 437 -204 438 -203
rect 438 -204 439 -203
rect 439 -204 440 -203
rect 440 -204 441 -203
rect 441 -204 442 -203
rect 442 -204 443 -203
rect 443 -204 444 -203
rect 444 -204 445 -203
rect 445 -204 446 -203
rect 446 -204 447 -203
rect 447 -204 448 -203
rect 448 -204 449 -203
rect 449 -204 450 -203
rect 450 -204 451 -203
rect 451 -204 452 -203
rect 452 -204 453 -203
rect 453 -204 454 -203
rect 454 -204 455 -203
rect 455 -204 456 -203
rect 456 -204 457 -203
rect 457 -204 458 -203
rect 458 -204 459 -203
rect 459 -204 460 -203
rect 460 -204 461 -203
rect 461 -204 462 -203
rect 462 -204 463 -203
rect 463 -204 464 -203
rect 464 -204 465 -203
rect 465 -204 466 -203
rect 466 -204 467 -203
rect 467 -204 468 -203
rect 468 -204 469 -203
rect 469 -204 470 -203
rect 470 -204 471 -203
rect 471 -204 472 -203
rect 472 -204 473 -203
rect 473 -204 474 -203
rect 474 -204 475 -203
rect 475 -204 476 -203
rect 476 -204 477 -203
rect 477 -204 478 -203
rect 478 -204 479 -203
rect 479 -204 480 -203
rect 2 -205 3 -204
rect 3 -205 4 -204
rect 4 -205 5 -204
rect 5 -205 6 -204
rect 6 -205 7 -204
rect 7 -205 8 -204
rect 8 -205 9 -204
rect 9 -205 10 -204
rect 10 -205 11 -204
rect 11 -205 12 -204
rect 12 -205 13 -204
rect 13 -205 14 -204
rect 14 -205 15 -204
rect 15 -205 16 -204
rect 16 -205 17 -204
rect 17 -205 18 -204
rect 18 -205 19 -204
rect 19 -205 20 -204
rect 20 -205 21 -204
rect 21 -205 22 -204
rect 22 -205 23 -204
rect 23 -205 24 -204
rect 24 -205 25 -204
rect 25 -205 26 -204
rect 26 -205 27 -204
rect 27 -205 28 -204
rect 28 -205 29 -204
rect 29 -205 30 -204
rect 30 -205 31 -204
rect 31 -205 32 -204
rect 32 -205 33 -204
rect 33 -205 34 -204
rect 34 -205 35 -204
rect 35 -205 36 -204
rect 36 -205 37 -204
rect 37 -205 38 -204
rect 38 -205 39 -204
rect 39 -205 40 -204
rect 40 -205 41 -204
rect 41 -205 42 -204
rect 42 -205 43 -204
rect 43 -205 44 -204
rect 44 -205 45 -204
rect 45 -205 46 -204
rect 46 -205 47 -204
rect 47 -205 48 -204
rect 48 -205 49 -204
rect 49 -205 50 -204
rect 50 -205 51 -204
rect 51 -205 52 -204
rect 52 -205 53 -204
rect 53 -205 54 -204
rect 54 -205 55 -204
rect 55 -205 56 -204
rect 56 -205 57 -204
rect 57 -205 58 -204
rect 58 -205 59 -204
rect 59 -205 60 -204
rect 60 -205 61 -204
rect 61 -205 62 -204
rect 62 -205 63 -204
rect 63 -205 64 -204
rect 64 -205 65 -204
rect 65 -205 66 -204
rect 66 -205 67 -204
rect 67 -205 68 -204
rect 68 -205 69 -204
rect 69 -205 70 -204
rect 70 -205 71 -204
rect 71 -205 72 -204
rect 72 -205 73 -204
rect 73 -205 74 -204
rect 74 -205 75 -204
rect 75 -205 76 -204
rect 76 -205 77 -204
rect 77 -205 78 -204
rect 78 -205 79 -204
rect 79 -205 80 -204
rect 80 -205 81 -204
rect 81 -205 82 -204
rect 82 -205 83 -204
rect 83 -205 84 -204
rect 84 -205 85 -204
rect 85 -205 86 -204
rect 86 -205 87 -204
rect 87 -205 88 -204
rect 88 -205 89 -204
rect 89 -205 90 -204
rect 90 -205 91 -204
rect 91 -205 92 -204
rect 92 -205 93 -204
rect 93 -205 94 -204
rect 94 -205 95 -204
rect 95 -205 96 -204
rect 96 -205 97 -204
rect 97 -205 98 -204
rect 98 -205 99 -204
rect 99 -205 100 -204
rect 100 -205 101 -204
rect 101 -205 102 -204
rect 102 -205 103 -204
rect 103 -205 104 -204
rect 104 -205 105 -204
rect 105 -205 106 -204
rect 106 -205 107 -204
rect 107 -205 108 -204
rect 108 -205 109 -204
rect 109 -205 110 -204
rect 110 -205 111 -204
rect 111 -205 112 -204
rect 112 -205 113 -204
rect 113 -205 114 -204
rect 114 -205 115 -204
rect 115 -205 116 -204
rect 116 -205 117 -204
rect 117 -205 118 -204
rect 118 -205 119 -204
rect 119 -205 120 -204
rect 120 -205 121 -204
rect 121 -205 122 -204
rect 122 -205 123 -204
rect 123 -205 124 -204
rect 124 -205 125 -204
rect 125 -205 126 -204
rect 126 -205 127 -204
rect 127 -205 128 -204
rect 128 -205 129 -204
rect 129 -205 130 -204
rect 130 -205 131 -204
rect 131 -205 132 -204
rect 132 -205 133 -204
rect 133 -205 134 -204
rect 134 -205 135 -204
rect 135 -205 136 -204
rect 136 -205 137 -204
rect 137 -205 138 -204
rect 138 -205 139 -204
rect 139 -205 140 -204
rect 140 -205 141 -204
rect 141 -205 142 -204
rect 142 -205 143 -204
rect 143 -205 144 -204
rect 144 -205 145 -204
rect 145 -205 146 -204
rect 146 -205 147 -204
rect 147 -205 148 -204
rect 148 -205 149 -204
rect 149 -205 150 -204
rect 150 -205 151 -204
rect 151 -205 152 -204
rect 152 -205 153 -204
rect 153 -205 154 -204
rect 154 -205 155 -204
rect 155 -205 156 -204
rect 156 -205 157 -204
rect 157 -205 158 -204
rect 158 -205 159 -204
rect 159 -205 160 -204
rect 160 -205 161 -204
rect 161 -205 162 -204
rect 162 -205 163 -204
rect 163 -205 164 -204
rect 164 -205 165 -204
rect 165 -205 166 -204
rect 166 -205 167 -204
rect 167 -205 168 -204
rect 168 -205 169 -204
rect 169 -205 170 -204
rect 170 -205 171 -204
rect 171 -205 172 -204
rect 172 -205 173 -204
rect 173 -205 174 -204
rect 174 -205 175 -204
rect 175 -205 176 -204
rect 176 -205 177 -204
rect 177 -205 178 -204
rect 178 -205 179 -204
rect 179 -205 180 -204
rect 180 -205 181 -204
rect 181 -205 182 -204
rect 182 -205 183 -204
rect 183 -205 184 -204
rect 184 -205 185 -204
rect 185 -205 186 -204
rect 186 -205 187 -204
rect 187 -205 188 -204
rect 188 -205 189 -204
rect 189 -205 190 -204
rect 190 -205 191 -204
rect 191 -205 192 -204
rect 192 -205 193 -204
rect 193 -205 194 -204
rect 194 -205 195 -204
rect 195 -205 196 -204
rect 196 -205 197 -204
rect 197 -205 198 -204
rect 198 -205 199 -204
rect 199 -205 200 -204
rect 200 -205 201 -204
rect 201 -205 202 -204
rect 202 -205 203 -204
rect 203 -205 204 -204
rect 204 -205 205 -204
rect 205 -205 206 -204
rect 206 -205 207 -204
rect 207 -205 208 -204
rect 208 -205 209 -204
rect 209 -205 210 -204
rect 210 -205 211 -204
rect 211 -205 212 -204
rect 212 -205 213 -204
rect 213 -205 214 -204
rect 214 -205 215 -204
rect 215 -205 216 -204
rect 216 -205 217 -204
rect 217 -205 218 -204
rect 218 -205 219 -204
rect 219 -205 220 -204
rect 220 -205 221 -204
rect 221 -205 222 -204
rect 222 -205 223 -204
rect 223 -205 224 -204
rect 224 -205 225 -204
rect 225 -205 226 -204
rect 226 -205 227 -204
rect 227 -205 228 -204
rect 228 -205 229 -204
rect 229 -205 230 -204
rect 230 -205 231 -204
rect 231 -205 232 -204
rect 232 -205 233 -204
rect 233 -205 234 -204
rect 234 -205 235 -204
rect 235 -205 236 -204
rect 236 -205 237 -204
rect 237 -205 238 -204
rect 238 -205 239 -204
rect 239 -205 240 -204
rect 240 -205 241 -204
rect 241 -205 242 -204
rect 242 -205 243 -204
rect 243 -205 244 -204
rect 244 -205 245 -204
rect 245 -205 246 -204
rect 246 -205 247 -204
rect 247 -205 248 -204
rect 248 -205 249 -204
rect 249 -205 250 -204
rect 250 -205 251 -204
rect 251 -205 252 -204
rect 252 -205 253 -204
rect 253 -205 254 -204
rect 254 -205 255 -204
rect 255 -205 256 -204
rect 256 -205 257 -204
rect 257 -205 258 -204
rect 258 -205 259 -204
rect 259 -205 260 -204
rect 260 -205 261 -204
rect 261 -205 262 -204
rect 262 -205 263 -204
rect 263 -205 264 -204
rect 264 -205 265 -204
rect 265 -205 266 -204
rect 266 -205 267 -204
rect 267 -205 268 -204
rect 268 -205 269 -204
rect 269 -205 270 -204
rect 270 -205 271 -204
rect 271 -205 272 -204
rect 272 -205 273 -204
rect 273 -205 274 -204
rect 274 -205 275 -204
rect 275 -205 276 -204
rect 276 -205 277 -204
rect 277 -205 278 -204
rect 278 -205 279 -204
rect 279 -205 280 -204
rect 280 -205 281 -204
rect 281 -205 282 -204
rect 282 -205 283 -204
rect 283 -205 284 -204
rect 284 -205 285 -204
rect 285 -205 286 -204
rect 286 -205 287 -204
rect 287 -205 288 -204
rect 288 -205 289 -204
rect 289 -205 290 -204
rect 290 -205 291 -204
rect 291 -205 292 -204
rect 292 -205 293 -204
rect 293 -205 294 -204
rect 294 -205 295 -204
rect 295 -205 296 -204
rect 296 -205 297 -204
rect 297 -205 298 -204
rect 298 -205 299 -204
rect 299 -205 300 -204
rect 300 -205 301 -204
rect 301 -205 302 -204
rect 302 -205 303 -204
rect 303 -205 304 -204
rect 304 -205 305 -204
rect 305 -205 306 -204
rect 306 -205 307 -204
rect 307 -205 308 -204
rect 308 -205 309 -204
rect 309 -205 310 -204
rect 310 -205 311 -204
rect 311 -205 312 -204
rect 312 -205 313 -204
rect 313 -205 314 -204
rect 314 -205 315 -204
rect 315 -205 316 -204
rect 316 -205 317 -204
rect 317 -205 318 -204
rect 318 -205 319 -204
rect 319 -205 320 -204
rect 320 -205 321 -204
rect 321 -205 322 -204
rect 322 -205 323 -204
rect 323 -205 324 -204
rect 324 -205 325 -204
rect 325 -205 326 -204
rect 326 -205 327 -204
rect 327 -205 328 -204
rect 328 -205 329 -204
rect 329 -205 330 -204
rect 330 -205 331 -204
rect 331 -205 332 -204
rect 332 -205 333 -204
rect 333 -205 334 -204
rect 334 -205 335 -204
rect 335 -205 336 -204
rect 336 -205 337 -204
rect 337 -205 338 -204
rect 338 -205 339 -204
rect 339 -205 340 -204
rect 340 -205 341 -204
rect 341 -205 342 -204
rect 342 -205 343 -204
rect 343 -205 344 -204
rect 344 -205 345 -204
rect 345 -205 346 -204
rect 346 -205 347 -204
rect 347 -205 348 -204
rect 348 -205 349 -204
rect 349 -205 350 -204
rect 350 -205 351 -204
rect 351 -205 352 -204
rect 352 -205 353 -204
rect 353 -205 354 -204
rect 354 -205 355 -204
rect 355 -205 356 -204
rect 356 -205 357 -204
rect 357 -205 358 -204
rect 358 -205 359 -204
rect 359 -205 360 -204
rect 360 -205 361 -204
rect 361 -205 362 -204
rect 362 -205 363 -204
rect 363 -205 364 -204
rect 364 -205 365 -204
rect 365 -205 366 -204
rect 366 -205 367 -204
rect 367 -205 368 -204
rect 368 -205 369 -204
rect 369 -205 370 -204
rect 370 -205 371 -204
rect 371 -205 372 -204
rect 372 -205 373 -204
rect 373 -205 374 -204
rect 374 -205 375 -204
rect 375 -205 376 -204
rect 376 -205 377 -204
rect 377 -205 378 -204
rect 378 -205 379 -204
rect 379 -205 380 -204
rect 380 -205 381 -204
rect 381 -205 382 -204
rect 382 -205 383 -204
rect 383 -205 384 -204
rect 384 -205 385 -204
rect 385 -205 386 -204
rect 386 -205 387 -204
rect 387 -205 388 -204
rect 388 -205 389 -204
rect 389 -205 390 -204
rect 390 -205 391 -204
rect 391 -205 392 -204
rect 392 -205 393 -204
rect 393 -205 394 -204
rect 394 -205 395 -204
rect 395 -205 396 -204
rect 396 -205 397 -204
rect 397 -205 398 -204
rect 398 -205 399 -204
rect 399 -205 400 -204
rect 400 -205 401 -204
rect 401 -205 402 -204
rect 402 -205 403 -204
rect 403 -205 404 -204
rect 404 -205 405 -204
rect 405 -205 406 -204
rect 406 -205 407 -204
rect 407 -205 408 -204
rect 408 -205 409 -204
rect 409 -205 410 -204
rect 410 -205 411 -204
rect 411 -205 412 -204
rect 412 -205 413 -204
rect 413 -205 414 -204
rect 414 -205 415 -204
rect 415 -205 416 -204
rect 416 -205 417 -204
rect 417 -205 418 -204
rect 418 -205 419 -204
rect 419 -205 420 -204
rect 420 -205 421 -204
rect 421 -205 422 -204
rect 422 -205 423 -204
rect 423 -205 424 -204
rect 424 -205 425 -204
rect 425 -205 426 -204
rect 426 -205 427 -204
rect 427 -205 428 -204
rect 428 -205 429 -204
rect 429 -205 430 -204
rect 430 -205 431 -204
rect 431 -205 432 -204
rect 432 -205 433 -204
rect 433 -205 434 -204
rect 434 -205 435 -204
rect 435 -205 436 -204
rect 436 -205 437 -204
rect 437 -205 438 -204
rect 438 -205 439 -204
rect 439 -205 440 -204
rect 440 -205 441 -204
rect 441 -205 442 -204
rect 442 -205 443 -204
rect 443 -205 444 -204
rect 444 -205 445 -204
rect 445 -205 446 -204
rect 446 -205 447 -204
rect 447 -205 448 -204
rect 448 -205 449 -204
rect 449 -205 450 -204
rect 450 -205 451 -204
rect 451 -205 452 -204
rect 452 -205 453 -204
rect 453 -205 454 -204
rect 454 -205 455 -204
rect 455 -205 456 -204
rect 456 -205 457 -204
rect 457 -205 458 -204
rect 458 -205 459 -204
rect 459 -205 460 -204
rect 460 -205 461 -204
rect 461 -205 462 -204
rect 462 -205 463 -204
rect 463 -205 464 -204
rect 464 -205 465 -204
rect 465 -205 466 -204
rect 466 -205 467 -204
rect 467 -205 468 -204
rect 468 -205 469 -204
rect 469 -205 470 -204
rect 470 -205 471 -204
rect 471 -205 472 -204
rect 472 -205 473 -204
rect 473 -205 474 -204
rect 474 -205 475 -204
rect 475 -205 476 -204
rect 476 -205 477 -204
rect 477 -205 478 -204
rect 478 -205 479 -204
rect 479 -205 480 -204
rect 2 -206 3 -205
rect 3 -206 4 -205
rect 4 -206 5 -205
rect 5 -206 6 -205
rect 6 -206 7 -205
rect 7 -206 8 -205
rect 8 -206 9 -205
rect 9 -206 10 -205
rect 10 -206 11 -205
rect 11 -206 12 -205
rect 12 -206 13 -205
rect 13 -206 14 -205
rect 14 -206 15 -205
rect 15 -206 16 -205
rect 16 -206 17 -205
rect 17 -206 18 -205
rect 18 -206 19 -205
rect 19 -206 20 -205
rect 20 -206 21 -205
rect 21 -206 22 -205
rect 22 -206 23 -205
rect 23 -206 24 -205
rect 24 -206 25 -205
rect 25 -206 26 -205
rect 26 -206 27 -205
rect 27 -206 28 -205
rect 28 -206 29 -205
rect 29 -206 30 -205
rect 30 -206 31 -205
rect 31 -206 32 -205
rect 32 -206 33 -205
rect 33 -206 34 -205
rect 34 -206 35 -205
rect 35 -206 36 -205
rect 36 -206 37 -205
rect 37 -206 38 -205
rect 38 -206 39 -205
rect 39 -206 40 -205
rect 40 -206 41 -205
rect 41 -206 42 -205
rect 42 -206 43 -205
rect 43 -206 44 -205
rect 44 -206 45 -205
rect 45 -206 46 -205
rect 46 -206 47 -205
rect 47 -206 48 -205
rect 48 -206 49 -205
rect 49 -206 50 -205
rect 50 -206 51 -205
rect 51 -206 52 -205
rect 52 -206 53 -205
rect 53 -206 54 -205
rect 54 -206 55 -205
rect 55 -206 56 -205
rect 56 -206 57 -205
rect 57 -206 58 -205
rect 58 -206 59 -205
rect 59 -206 60 -205
rect 60 -206 61 -205
rect 61 -206 62 -205
rect 62 -206 63 -205
rect 63 -206 64 -205
rect 64 -206 65 -205
rect 65 -206 66 -205
rect 66 -206 67 -205
rect 67 -206 68 -205
rect 68 -206 69 -205
rect 69 -206 70 -205
rect 70 -206 71 -205
rect 71 -206 72 -205
rect 72 -206 73 -205
rect 73 -206 74 -205
rect 74 -206 75 -205
rect 75 -206 76 -205
rect 76 -206 77 -205
rect 77 -206 78 -205
rect 78 -206 79 -205
rect 79 -206 80 -205
rect 80 -206 81 -205
rect 81 -206 82 -205
rect 82 -206 83 -205
rect 83 -206 84 -205
rect 84 -206 85 -205
rect 85 -206 86 -205
rect 86 -206 87 -205
rect 87 -206 88 -205
rect 88 -206 89 -205
rect 89 -206 90 -205
rect 90 -206 91 -205
rect 91 -206 92 -205
rect 92 -206 93 -205
rect 93 -206 94 -205
rect 94 -206 95 -205
rect 95 -206 96 -205
rect 96 -206 97 -205
rect 97 -206 98 -205
rect 98 -206 99 -205
rect 99 -206 100 -205
rect 100 -206 101 -205
rect 101 -206 102 -205
rect 102 -206 103 -205
rect 103 -206 104 -205
rect 104 -206 105 -205
rect 105 -206 106 -205
rect 106 -206 107 -205
rect 107 -206 108 -205
rect 108 -206 109 -205
rect 109 -206 110 -205
rect 110 -206 111 -205
rect 111 -206 112 -205
rect 112 -206 113 -205
rect 113 -206 114 -205
rect 114 -206 115 -205
rect 115 -206 116 -205
rect 116 -206 117 -205
rect 117 -206 118 -205
rect 118 -206 119 -205
rect 119 -206 120 -205
rect 120 -206 121 -205
rect 121 -206 122 -205
rect 122 -206 123 -205
rect 123 -206 124 -205
rect 124 -206 125 -205
rect 125 -206 126 -205
rect 126 -206 127 -205
rect 127 -206 128 -205
rect 128 -206 129 -205
rect 129 -206 130 -205
rect 130 -206 131 -205
rect 131 -206 132 -205
rect 132 -206 133 -205
rect 133 -206 134 -205
rect 134 -206 135 -205
rect 135 -206 136 -205
rect 136 -206 137 -205
rect 137 -206 138 -205
rect 138 -206 139 -205
rect 139 -206 140 -205
rect 140 -206 141 -205
rect 141 -206 142 -205
rect 142 -206 143 -205
rect 143 -206 144 -205
rect 144 -206 145 -205
rect 145 -206 146 -205
rect 146 -206 147 -205
rect 147 -206 148 -205
rect 148 -206 149 -205
rect 149 -206 150 -205
rect 150 -206 151 -205
rect 151 -206 152 -205
rect 152 -206 153 -205
rect 153 -206 154 -205
rect 154 -206 155 -205
rect 155 -206 156 -205
rect 156 -206 157 -205
rect 157 -206 158 -205
rect 158 -206 159 -205
rect 159 -206 160 -205
rect 160 -206 161 -205
rect 161 -206 162 -205
rect 162 -206 163 -205
rect 163 -206 164 -205
rect 164 -206 165 -205
rect 165 -206 166 -205
rect 166 -206 167 -205
rect 167 -206 168 -205
rect 168 -206 169 -205
rect 169 -206 170 -205
rect 170 -206 171 -205
rect 171 -206 172 -205
rect 172 -206 173 -205
rect 173 -206 174 -205
rect 174 -206 175 -205
rect 175 -206 176 -205
rect 176 -206 177 -205
rect 177 -206 178 -205
rect 178 -206 179 -205
rect 179 -206 180 -205
rect 180 -206 181 -205
rect 181 -206 182 -205
rect 182 -206 183 -205
rect 183 -206 184 -205
rect 184 -206 185 -205
rect 185 -206 186 -205
rect 186 -206 187 -205
rect 187 -206 188 -205
rect 188 -206 189 -205
rect 189 -206 190 -205
rect 190 -206 191 -205
rect 191 -206 192 -205
rect 192 -206 193 -205
rect 193 -206 194 -205
rect 194 -206 195 -205
rect 195 -206 196 -205
rect 196 -206 197 -205
rect 197 -206 198 -205
rect 198 -206 199 -205
rect 199 -206 200 -205
rect 200 -206 201 -205
rect 201 -206 202 -205
rect 202 -206 203 -205
rect 203 -206 204 -205
rect 204 -206 205 -205
rect 205 -206 206 -205
rect 206 -206 207 -205
rect 207 -206 208 -205
rect 208 -206 209 -205
rect 209 -206 210 -205
rect 210 -206 211 -205
rect 211 -206 212 -205
rect 212 -206 213 -205
rect 213 -206 214 -205
rect 214 -206 215 -205
rect 215 -206 216 -205
rect 216 -206 217 -205
rect 217 -206 218 -205
rect 218 -206 219 -205
rect 219 -206 220 -205
rect 220 -206 221 -205
rect 221 -206 222 -205
rect 222 -206 223 -205
rect 223 -206 224 -205
rect 224 -206 225 -205
rect 225 -206 226 -205
rect 226 -206 227 -205
rect 227 -206 228 -205
rect 228 -206 229 -205
rect 229 -206 230 -205
rect 230 -206 231 -205
rect 231 -206 232 -205
rect 232 -206 233 -205
rect 233 -206 234 -205
rect 234 -206 235 -205
rect 235 -206 236 -205
rect 236 -206 237 -205
rect 237 -206 238 -205
rect 238 -206 239 -205
rect 239 -206 240 -205
rect 240 -206 241 -205
rect 241 -206 242 -205
rect 242 -206 243 -205
rect 243 -206 244 -205
rect 244 -206 245 -205
rect 245 -206 246 -205
rect 246 -206 247 -205
rect 247 -206 248 -205
rect 248 -206 249 -205
rect 249 -206 250 -205
rect 250 -206 251 -205
rect 251 -206 252 -205
rect 252 -206 253 -205
rect 253 -206 254 -205
rect 254 -206 255 -205
rect 255 -206 256 -205
rect 256 -206 257 -205
rect 257 -206 258 -205
rect 258 -206 259 -205
rect 259 -206 260 -205
rect 260 -206 261 -205
rect 261 -206 262 -205
rect 262 -206 263 -205
rect 263 -206 264 -205
rect 264 -206 265 -205
rect 265 -206 266 -205
rect 266 -206 267 -205
rect 267 -206 268 -205
rect 268 -206 269 -205
rect 269 -206 270 -205
rect 270 -206 271 -205
rect 271 -206 272 -205
rect 272 -206 273 -205
rect 273 -206 274 -205
rect 274 -206 275 -205
rect 275 -206 276 -205
rect 276 -206 277 -205
rect 277 -206 278 -205
rect 278 -206 279 -205
rect 279 -206 280 -205
rect 280 -206 281 -205
rect 281 -206 282 -205
rect 282 -206 283 -205
rect 283 -206 284 -205
rect 284 -206 285 -205
rect 285 -206 286 -205
rect 286 -206 287 -205
rect 287 -206 288 -205
rect 288 -206 289 -205
rect 289 -206 290 -205
rect 290 -206 291 -205
rect 291 -206 292 -205
rect 292 -206 293 -205
rect 293 -206 294 -205
rect 294 -206 295 -205
rect 295 -206 296 -205
rect 296 -206 297 -205
rect 297 -206 298 -205
rect 298 -206 299 -205
rect 299 -206 300 -205
rect 300 -206 301 -205
rect 301 -206 302 -205
rect 302 -206 303 -205
rect 303 -206 304 -205
rect 304 -206 305 -205
rect 305 -206 306 -205
rect 306 -206 307 -205
rect 307 -206 308 -205
rect 308 -206 309 -205
rect 309 -206 310 -205
rect 310 -206 311 -205
rect 311 -206 312 -205
rect 312 -206 313 -205
rect 313 -206 314 -205
rect 314 -206 315 -205
rect 315 -206 316 -205
rect 316 -206 317 -205
rect 317 -206 318 -205
rect 318 -206 319 -205
rect 319 -206 320 -205
rect 320 -206 321 -205
rect 321 -206 322 -205
rect 322 -206 323 -205
rect 323 -206 324 -205
rect 324 -206 325 -205
rect 325 -206 326 -205
rect 326 -206 327 -205
rect 327 -206 328 -205
rect 328 -206 329 -205
rect 329 -206 330 -205
rect 330 -206 331 -205
rect 331 -206 332 -205
rect 332 -206 333 -205
rect 333 -206 334 -205
rect 334 -206 335 -205
rect 335 -206 336 -205
rect 336 -206 337 -205
rect 337 -206 338 -205
rect 338 -206 339 -205
rect 339 -206 340 -205
rect 340 -206 341 -205
rect 341 -206 342 -205
rect 342 -206 343 -205
rect 343 -206 344 -205
rect 344 -206 345 -205
rect 345 -206 346 -205
rect 346 -206 347 -205
rect 347 -206 348 -205
rect 348 -206 349 -205
rect 349 -206 350 -205
rect 350 -206 351 -205
rect 351 -206 352 -205
rect 352 -206 353 -205
rect 353 -206 354 -205
rect 354 -206 355 -205
rect 355 -206 356 -205
rect 356 -206 357 -205
rect 357 -206 358 -205
rect 358 -206 359 -205
rect 359 -206 360 -205
rect 360 -206 361 -205
rect 361 -206 362 -205
rect 362 -206 363 -205
rect 363 -206 364 -205
rect 364 -206 365 -205
rect 365 -206 366 -205
rect 366 -206 367 -205
rect 367 -206 368 -205
rect 368 -206 369 -205
rect 369 -206 370 -205
rect 370 -206 371 -205
rect 371 -206 372 -205
rect 372 -206 373 -205
rect 373 -206 374 -205
rect 374 -206 375 -205
rect 375 -206 376 -205
rect 376 -206 377 -205
rect 377 -206 378 -205
rect 378 -206 379 -205
rect 379 -206 380 -205
rect 380 -206 381 -205
rect 381 -206 382 -205
rect 382 -206 383 -205
rect 383 -206 384 -205
rect 384 -206 385 -205
rect 385 -206 386 -205
rect 386 -206 387 -205
rect 387 -206 388 -205
rect 388 -206 389 -205
rect 389 -206 390 -205
rect 390 -206 391 -205
rect 391 -206 392 -205
rect 392 -206 393 -205
rect 393 -206 394 -205
rect 394 -206 395 -205
rect 395 -206 396 -205
rect 396 -206 397 -205
rect 397 -206 398 -205
rect 398 -206 399 -205
rect 399 -206 400 -205
rect 400 -206 401 -205
rect 401 -206 402 -205
rect 402 -206 403 -205
rect 403 -206 404 -205
rect 404 -206 405 -205
rect 405 -206 406 -205
rect 406 -206 407 -205
rect 407 -206 408 -205
rect 408 -206 409 -205
rect 409 -206 410 -205
rect 410 -206 411 -205
rect 411 -206 412 -205
rect 412 -206 413 -205
rect 413 -206 414 -205
rect 414 -206 415 -205
rect 415 -206 416 -205
rect 416 -206 417 -205
rect 417 -206 418 -205
rect 418 -206 419 -205
rect 419 -206 420 -205
rect 420 -206 421 -205
rect 421 -206 422 -205
rect 422 -206 423 -205
rect 423 -206 424 -205
rect 424 -206 425 -205
rect 425 -206 426 -205
rect 426 -206 427 -205
rect 427 -206 428 -205
rect 428 -206 429 -205
rect 429 -206 430 -205
rect 430 -206 431 -205
rect 431 -206 432 -205
rect 432 -206 433 -205
rect 433 -206 434 -205
rect 434 -206 435 -205
rect 435 -206 436 -205
rect 436 -206 437 -205
rect 437 -206 438 -205
rect 438 -206 439 -205
rect 439 -206 440 -205
rect 440 -206 441 -205
rect 441 -206 442 -205
rect 442 -206 443 -205
rect 443 -206 444 -205
rect 444 -206 445 -205
rect 445 -206 446 -205
rect 446 -206 447 -205
rect 447 -206 448 -205
rect 448 -206 449 -205
rect 449 -206 450 -205
rect 450 -206 451 -205
rect 451 -206 452 -205
rect 452 -206 453 -205
rect 453 -206 454 -205
rect 454 -206 455 -205
rect 455 -206 456 -205
rect 456 -206 457 -205
rect 457 -206 458 -205
rect 458 -206 459 -205
rect 459 -206 460 -205
rect 460 -206 461 -205
rect 461 -206 462 -205
rect 462 -206 463 -205
rect 463 -206 464 -205
rect 464 -206 465 -205
rect 465 -206 466 -205
rect 466 -206 467 -205
rect 467 -206 468 -205
rect 468 -206 469 -205
rect 469 -206 470 -205
rect 470 -206 471 -205
rect 471 -206 472 -205
rect 472 -206 473 -205
rect 473 -206 474 -205
rect 474 -206 475 -205
rect 475 -206 476 -205
rect 476 -206 477 -205
rect 477 -206 478 -205
rect 478 -206 479 -205
rect 479 -206 480 -205
rect 2 -207 3 -206
rect 3 -207 4 -206
rect 4 -207 5 -206
rect 5 -207 6 -206
rect 6 -207 7 -206
rect 7 -207 8 -206
rect 8 -207 9 -206
rect 9 -207 10 -206
rect 10 -207 11 -206
rect 11 -207 12 -206
rect 12 -207 13 -206
rect 13 -207 14 -206
rect 14 -207 15 -206
rect 15 -207 16 -206
rect 16 -207 17 -206
rect 17 -207 18 -206
rect 18 -207 19 -206
rect 19 -207 20 -206
rect 20 -207 21 -206
rect 21 -207 22 -206
rect 22 -207 23 -206
rect 23 -207 24 -206
rect 24 -207 25 -206
rect 25 -207 26 -206
rect 26 -207 27 -206
rect 27 -207 28 -206
rect 28 -207 29 -206
rect 29 -207 30 -206
rect 30 -207 31 -206
rect 31 -207 32 -206
rect 32 -207 33 -206
rect 33 -207 34 -206
rect 34 -207 35 -206
rect 35 -207 36 -206
rect 36 -207 37 -206
rect 37 -207 38 -206
rect 38 -207 39 -206
rect 39 -207 40 -206
rect 40 -207 41 -206
rect 41 -207 42 -206
rect 42 -207 43 -206
rect 43 -207 44 -206
rect 44 -207 45 -206
rect 45 -207 46 -206
rect 46 -207 47 -206
rect 47 -207 48 -206
rect 48 -207 49 -206
rect 49 -207 50 -206
rect 50 -207 51 -206
rect 51 -207 52 -206
rect 52 -207 53 -206
rect 53 -207 54 -206
rect 54 -207 55 -206
rect 55 -207 56 -206
rect 56 -207 57 -206
rect 57 -207 58 -206
rect 58 -207 59 -206
rect 59 -207 60 -206
rect 60 -207 61 -206
rect 61 -207 62 -206
rect 62 -207 63 -206
rect 63 -207 64 -206
rect 64 -207 65 -206
rect 65 -207 66 -206
rect 66 -207 67 -206
rect 67 -207 68 -206
rect 68 -207 69 -206
rect 69 -207 70 -206
rect 70 -207 71 -206
rect 71 -207 72 -206
rect 72 -207 73 -206
rect 73 -207 74 -206
rect 74 -207 75 -206
rect 75 -207 76 -206
rect 76 -207 77 -206
rect 77 -207 78 -206
rect 78 -207 79 -206
rect 79 -207 80 -206
rect 80 -207 81 -206
rect 81 -207 82 -206
rect 82 -207 83 -206
rect 83 -207 84 -206
rect 84 -207 85 -206
rect 85 -207 86 -206
rect 86 -207 87 -206
rect 87 -207 88 -206
rect 88 -207 89 -206
rect 89 -207 90 -206
rect 90 -207 91 -206
rect 91 -207 92 -206
rect 92 -207 93 -206
rect 93 -207 94 -206
rect 94 -207 95 -206
rect 95 -207 96 -206
rect 96 -207 97 -206
rect 97 -207 98 -206
rect 98 -207 99 -206
rect 99 -207 100 -206
rect 100 -207 101 -206
rect 101 -207 102 -206
rect 102 -207 103 -206
rect 103 -207 104 -206
rect 104 -207 105 -206
rect 105 -207 106 -206
rect 106 -207 107 -206
rect 107 -207 108 -206
rect 108 -207 109 -206
rect 109 -207 110 -206
rect 110 -207 111 -206
rect 111 -207 112 -206
rect 112 -207 113 -206
rect 113 -207 114 -206
rect 114 -207 115 -206
rect 115 -207 116 -206
rect 116 -207 117 -206
rect 117 -207 118 -206
rect 118 -207 119 -206
rect 119 -207 120 -206
rect 120 -207 121 -206
rect 121 -207 122 -206
rect 122 -207 123 -206
rect 123 -207 124 -206
rect 124 -207 125 -206
rect 125 -207 126 -206
rect 126 -207 127 -206
rect 127 -207 128 -206
rect 128 -207 129 -206
rect 129 -207 130 -206
rect 130 -207 131 -206
rect 131 -207 132 -206
rect 132 -207 133 -206
rect 133 -207 134 -206
rect 134 -207 135 -206
rect 135 -207 136 -206
rect 136 -207 137 -206
rect 137 -207 138 -206
rect 138 -207 139 -206
rect 139 -207 140 -206
rect 140 -207 141 -206
rect 141 -207 142 -206
rect 142 -207 143 -206
rect 143 -207 144 -206
rect 144 -207 145 -206
rect 145 -207 146 -206
rect 146 -207 147 -206
rect 147 -207 148 -206
rect 148 -207 149 -206
rect 149 -207 150 -206
rect 150 -207 151 -206
rect 151 -207 152 -206
rect 152 -207 153 -206
rect 153 -207 154 -206
rect 154 -207 155 -206
rect 155 -207 156 -206
rect 156 -207 157 -206
rect 157 -207 158 -206
rect 158 -207 159 -206
rect 159 -207 160 -206
rect 160 -207 161 -206
rect 161 -207 162 -206
rect 162 -207 163 -206
rect 163 -207 164 -206
rect 164 -207 165 -206
rect 165 -207 166 -206
rect 166 -207 167 -206
rect 167 -207 168 -206
rect 168 -207 169 -206
rect 169 -207 170 -206
rect 170 -207 171 -206
rect 171 -207 172 -206
rect 172 -207 173 -206
rect 173 -207 174 -206
rect 174 -207 175 -206
rect 175 -207 176 -206
rect 176 -207 177 -206
rect 177 -207 178 -206
rect 178 -207 179 -206
rect 179 -207 180 -206
rect 180 -207 181 -206
rect 181 -207 182 -206
rect 182 -207 183 -206
rect 183 -207 184 -206
rect 184 -207 185 -206
rect 185 -207 186 -206
rect 186 -207 187 -206
rect 187 -207 188 -206
rect 188 -207 189 -206
rect 189 -207 190 -206
rect 190 -207 191 -206
rect 191 -207 192 -206
rect 192 -207 193 -206
rect 193 -207 194 -206
rect 194 -207 195 -206
rect 195 -207 196 -206
rect 196 -207 197 -206
rect 197 -207 198 -206
rect 198 -207 199 -206
rect 199 -207 200 -206
rect 200 -207 201 -206
rect 201 -207 202 -206
rect 202 -207 203 -206
rect 203 -207 204 -206
rect 204 -207 205 -206
rect 205 -207 206 -206
rect 206 -207 207 -206
rect 207 -207 208 -206
rect 208 -207 209 -206
rect 209 -207 210 -206
rect 210 -207 211 -206
rect 211 -207 212 -206
rect 212 -207 213 -206
rect 213 -207 214 -206
rect 214 -207 215 -206
rect 215 -207 216 -206
rect 216 -207 217 -206
rect 217 -207 218 -206
rect 218 -207 219 -206
rect 219 -207 220 -206
rect 220 -207 221 -206
rect 221 -207 222 -206
rect 222 -207 223 -206
rect 223 -207 224 -206
rect 224 -207 225 -206
rect 225 -207 226 -206
rect 226 -207 227 -206
rect 227 -207 228 -206
rect 228 -207 229 -206
rect 229 -207 230 -206
rect 230 -207 231 -206
rect 231 -207 232 -206
rect 232 -207 233 -206
rect 233 -207 234 -206
rect 234 -207 235 -206
rect 235 -207 236 -206
rect 236 -207 237 -206
rect 237 -207 238 -206
rect 238 -207 239 -206
rect 239 -207 240 -206
rect 240 -207 241 -206
rect 241 -207 242 -206
rect 242 -207 243 -206
rect 243 -207 244 -206
rect 244 -207 245 -206
rect 245 -207 246 -206
rect 246 -207 247 -206
rect 247 -207 248 -206
rect 248 -207 249 -206
rect 249 -207 250 -206
rect 250 -207 251 -206
rect 251 -207 252 -206
rect 252 -207 253 -206
rect 253 -207 254 -206
rect 254 -207 255 -206
rect 255 -207 256 -206
rect 256 -207 257 -206
rect 257 -207 258 -206
rect 258 -207 259 -206
rect 259 -207 260 -206
rect 260 -207 261 -206
rect 261 -207 262 -206
rect 262 -207 263 -206
rect 263 -207 264 -206
rect 264 -207 265 -206
rect 265 -207 266 -206
rect 266 -207 267 -206
rect 267 -207 268 -206
rect 268 -207 269 -206
rect 269 -207 270 -206
rect 270 -207 271 -206
rect 271 -207 272 -206
rect 272 -207 273 -206
rect 273 -207 274 -206
rect 274 -207 275 -206
rect 275 -207 276 -206
rect 276 -207 277 -206
rect 277 -207 278 -206
rect 278 -207 279 -206
rect 279 -207 280 -206
rect 280 -207 281 -206
rect 281 -207 282 -206
rect 282 -207 283 -206
rect 283 -207 284 -206
rect 284 -207 285 -206
rect 285 -207 286 -206
rect 286 -207 287 -206
rect 287 -207 288 -206
rect 288 -207 289 -206
rect 289 -207 290 -206
rect 290 -207 291 -206
rect 291 -207 292 -206
rect 292 -207 293 -206
rect 293 -207 294 -206
rect 294 -207 295 -206
rect 295 -207 296 -206
rect 296 -207 297 -206
rect 297 -207 298 -206
rect 298 -207 299 -206
rect 299 -207 300 -206
rect 300 -207 301 -206
rect 301 -207 302 -206
rect 302 -207 303 -206
rect 303 -207 304 -206
rect 304 -207 305 -206
rect 305 -207 306 -206
rect 306 -207 307 -206
rect 307 -207 308 -206
rect 308 -207 309 -206
rect 309 -207 310 -206
rect 310 -207 311 -206
rect 311 -207 312 -206
rect 312 -207 313 -206
rect 313 -207 314 -206
rect 314 -207 315 -206
rect 315 -207 316 -206
rect 316 -207 317 -206
rect 317 -207 318 -206
rect 318 -207 319 -206
rect 319 -207 320 -206
rect 320 -207 321 -206
rect 321 -207 322 -206
rect 322 -207 323 -206
rect 323 -207 324 -206
rect 324 -207 325 -206
rect 325 -207 326 -206
rect 326 -207 327 -206
rect 327 -207 328 -206
rect 328 -207 329 -206
rect 329 -207 330 -206
rect 330 -207 331 -206
rect 331 -207 332 -206
rect 332 -207 333 -206
rect 333 -207 334 -206
rect 334 -207 335 -206
rect 335 -207 336 -206
rect 336 -207 337 -206
rect 337 -207 338 -206
rect 338 -207 339 -206
rect 339 -207 340 -206
rect 340 -207 341 -206
rect 341 -207 342 -206
rect 342 -207 343 -206
rect 343 -207 344 -206
rect 344 -207 345 -206
rect 345 -207 346 -206
rect 346 -207 347 -206
rect 347 -207 348 -206
rect 348 -207 349 -206
rect 349 -207 350 -206
rect 350 -207 351 -206
rect 351 -207 352 -206
rect 352 -207 353 -206
rect 353 -207 354 -206
rect 354 -207 355 -206
rect 355 -207 356 -206
rect 356 -207 357 -206
rect 357 -207 358 -206
rect 358 -207 359 -206
rect 359 -207 360 -206
rect 360 -207 361 -206
rect 361 -207 362 -206
rect 362 -207 363 -206
rect 363 -207 364 -206
rect 364 -207 365 -206
rect 365 -207 366 -206
rect 366 -207 367 -206
rect 367 -207 368 -206
rect 368 -207 369 -206
rect 369 -207 370 -206
rect 370 -207 371 -206
rect 371 -207 372 -206
rect 372 -207 373 -206
rect 373 -207 374 -206
rect 374 -207 375 -206
rect 375 -207 376 -206
rect 376 -207 377 -206
rect 377 -207 378 -206
rect 378 -207 379 -206
rect 379 -207 380 -206
rect 380 -207 381 -206
rect 381 -207 382 -206
rect 382 -207 383 -206
rect 383 -207 384 -206
rect 384 -207 385 -206
rect 385 -207 386 -206
rect 386 -207 387 -206
rect 387 -207 388 -206
rect 388 -207 389 -206
rect 389 -207 390 -206
rect 390 -207 391 -206
rect 391 -207 392 -206
rect 392 -207 393 -206
rect 393 -207 394 -206
rect 394 -207 395 -206
rect 395 -207 396 -206
rect 396 -207 397 -206
rect 397 -207 398 -206
rect 398 -207 399 -206
rect 399 -207 400 -206
rect 400 -207 401 -206
rect 401 -207 402 -206
rect 402 -207 403 -206
rect 403 -207 404 -206
rect 404 -207 405 -206
rect 405 -207 406 -206
rect 406 -207 407 -206
rect 407 -207 408 -206
rect 408 -207 409 -206
rect 409 -207 410 -206
rect 410 -207 411 -206
rect 411 -207 412 -206
rect 412 -207 413 -206
rect 413 -207 414 -206
rect 414 -207 415 -206
rect 415 -207 416 -206
rect 416 -207 417 -206
rect 417 -207 418 -206
rect 418 -207 419 -206
rect 419 -207 420 -206
rect 420 -207 421 -206
rect 421 -207 422 -206
rect 422 -207 423 -206
rect 423 -207 424 -206
rect 424 -207 425 -206
rect 425 -207 426 -206
rect 426 -207 427 -206
rect 427 -207 428 -206
rect 428 -207 429 -206
rect 429 -207 430 -206
rect 430 -207 431 -206
rect 431 -207 432 -206
rect 432 -207 433 -206
rect 433 -207 434 -206
rect 434 -207 435 -206
rect 435 -207 436 -206
rect 436 -207 437 -206
rect 437 -207 438 -206
rect 438 -207 439 -206
rect 439 -207 440 -206
rect 440 -207 441 -206
rect 441 -207 442 -206
rect 442 -207 443 -206
rect 443 -207 444 -206
rect 444 -207 445 -206
rect 445 -207 446 -206
rect 446 -207 447 -206
rect 447 -207 448 -206
rect 448 -207 449 -206
rect 449 -207 450 -206
rect 450 -207 451 -206
rect 451 -207 452 -206
rect 452 -207 453 -206
rect 453 -207 454 -206
rect 454 -207 455 -206
rect 455 -207 456 -206
rect 456 -207 457 -206
rect 457 -207 458 -206
rect 458 -207 459 -206
rect 459 -207 460 -206
rect 460 -207 461 -206
rect 461 -207 462 -206
rect 462 -207 463 -206
rect 463 -207 464 -206
rect 464 -207 465 -206
rect 465 -207 466 -206
rect 466 -207 467 -206
rect 467 -207 468 -206
rect 468 -207 469 -206
rect 469 -207 470 -206
rect 470 -207 471 -206
rect 471 -207 472 -206
rect 472 -207 473 -206
rect 473 -207 474 -206
rect 474 -207 475 -206
rect 475 -207 476 -206
rect 476 -207 477 -206
rect 477 -207 478 -206
rect 478 -207 479 -206
rect 479 -207 480 -206
rect 2 -208 3 -207
rect 3 -208 4 -207
rect 4 -208 5 -207
rect 5 -208 6 -207
rect 6 -208 7 -207
rect 7 -208 8 -207
rect 8 -208 9 -207
rect 9 -208 10 -207
rect 10 -208 11 -207
rect 11 -208 12 -207
rect 12 -208 13 -207
rect 13 -208 14 -207
rect 14 -208 15 -207
rect 15 -208 16 -207
rect 16 -208 17 -207
rect 17 -208 18 -207
rect 18 -208 19 -207
rect 19 -208 20 -207
rect 20 -208 21 -207
rect 21 -208 22 -207
rect 22 -208 23 -207
rect 23 -208 24 -207
rect 24 -208 25 -207
rect 25 -208 26 -207
rect 26 -208 27 -207
rect 27 -208 28 -207
rect 28 -208 29 -207
rect 29 -208 30 -207
rect 30 -208 31 -207
rect 31 -208 32 -207
rect 32 -208 33 -207
rect 33 -208 34 -207
rect 34 -208 35 -207
rect 35 -208 36 -207
rect 36 -208 37 -207
rect 37 -208 38 -207
rect 38 -208 39 -207
rect 39 -208 40 -207
rect 40 -208 41 -207
rect 41 -208 42 -207
rect 42 -208 43 -207
rect 43 -208 44 -207
rect 44 -208 45 -207
rect 45 -208 46 -207
rect 46 -208 47 -207
rect 47 -208 48 -207
rect 48 -208 49 -207
rect 49 -208 50 -207
rect 50 -208 51 -207
rect 51 -208 52 -207
rect 52 -208 53 -207
rect 53 -208 54 -207
rect 54 -208 55 -207
rect 55 -208 56 -207
rect 56 -208 57 -207
rect 57 -208 58 -207
rect 58 -208 59 -207
rect 59 -208 60 -207
rect 60 -208 61 -207
rect 61 -208 62 -207
rect 62 -208 63 -207
rect 63 -208 64 -207
rect 64 -208 65 -207
rect 65 -208 66 -207
rect 66 -208 67 -207
rect 67 -208 68 -207
rect 68 -208 69 -207
rect 69 -208 70 -207
rect 70 -208 71 -207
rect 71 -208 72 -207
rect 72 -208 73 -207
rect 73 -208 74 -207
rect 74 -208 75 -207
rect 75 -208 76 -207
rect 76 -208 77 -207
rect 77 -208 78 -207
rect 78 -208 79 -207
rect 79 -208 80 -207
rect 80 -208 81 -207
rect 81 -208 82 -207
rect 82 -208 83 -207
rect 83 -208 84 -207
rect 84 -208 85 -207
rect 85 -208 86 -207
rect 86 -208 87 -207
rect 87 -208 88 -207
rect 88 -208 89 -207
rect 89 -208 90 -207
rect 90 -208 91 -207
rect 91 -208 92 -207
rect 92 -208 93 -207
rect 93 -208 94 -207
rect 94 -208 95 -207
rect 95 -208 96 -207
rect 96 -208 97 -207
rect 97 -208 98 -207
rect 98 -208 99 -207
rect 99 -208 100 -207
rect 100 -208 101 -207
rect 101 -208 102 -207
rect 102 -208 103 -207
rect 103 -208 104 -207
rect 104 -208 105 -207
rect 105 -208 106 -207
rect 106 -208 107 -207
rect 107 -208 108 -207
rect 108 -208 109 -207
rect 109 -208 110 -207
rect 110 -208 111 -207
rect 111 -208 112 -207
rect 112 -208 113 -207
rect 113 -208 114 -207
rect 114 -208 115 -207
rect 115 -208 116 -207
rect 116 -208 117 -207
rect 117 -208 118 -207
rect 118 -208 119 -207
rect 119 -208 120 -207
rect 120 -208 121 -207
rect 121 -208 122 -207
rect 122 -208 123 -207
rect 123 -208 124 -207
rect 124 -208 125 -207
rect 125 -208 126 -207
rect 126 -208 127 -207
rect 127 -208 128 -207
rect 128 -208 129 -207
rect 129 -208 130 -207
rect 130 -208 131 -207
rect 131 -208 132 -207
rect 132 -208 133 -207
rect 133 -208 134 -207
rect 134 -208 135 -207
rect 135 -208 136 -207
rect 136 -208 137 -207
rect 137 -208 138 -207
rect 138 -208 139 -207
rect 139 -208 140 -207
rect 140 -208 141 -207
rect 141 -208 142 -207
rect 142 -208 143 -207
rect 143 -208 144 -207
rect 144 -208 145 -207
rect 145 -208 146 -207
rect 146 -208 147 -207
rect 147 -208 148 -207
rect 148 -208 149 -207
rect 149 -208 150 -207
rect 150 -208 151 -207
rect 151 -208 152 -207
rect 152 -208 153 -207
rect 153 -208 154 -207
rect 154 -208 155 -207
rect 155 -208 156 -207
rect 156 -208 157 -207
rect 157 -208 158 -207
rect 158 -208 159 -207
rect 159 -208 160 -207
rect 160 -208 161 -207
rect 161 -208 162 -207
rect 162 -208 163 -207
rect 163 -208 164 -207
rect 164 -208 165 -207
rect 165 -208 166 -207
rect 166 -208 167 -207
rect 167 -208 168 -207
rect 168 -208 169 -207
rect 169 -208 170 -207
rect 170 -208 171 -207
rect 171 -208 172 -207
rect 172 -208 173 -207
rect 173 -208 174 -207
rect 174 -208 175 -207
rect 175 -208 176 -207
rect 176 -208 177 -207
rect 177 -208 178 -207
rect 178 -208 179 -207
rect 179 -208 180 -207
rect 180 -208 181 -207
rect 181 -208 182 -207
rect 182 -208 183 -207
rect 183 -208 184 -207
rect 184 -208 185 -207
rect 185 -208 186 -207
rect 186 -208 187 -207
rect 187 -208 188 -207
rect 188 -208 189 -207
rect 189 -208 190 -207
rect 190 -208 191 -207
rect 191 -208 192 -207
rect 192 -208 193 -207
rect 193 -208 194 -207
rect 194 -208 195 -207
rect 195 -208 196 -207
rect 196 -208 197 -207
rect 197 -208 198 -207
rect 198 -208 199 -207
rect 199 -208 200 -207
rect 200 -208 201 -207
rect 201 -208 202 -207
rect 202 -208 203 -207
rect 203 -208 204 -207
rect 204 -208 205 -207
rect 205 -208 206 -207
rect 206 -208 207 -207
rect 207 -208 208 -207
rect 208 -208 209 -207
rect 209 -208 210 -207
rect 210 -208 211 -207
rect 211 -208 212 -207
rect 212 -208 213 -207
rect 213 -208 214 -207
rect 214 -208 215 -207
rect 215 -208 216 -207
rect 216 -208 217 -207
rect 217 -208 218 -207
rect 218 -208 219 -207
rect 219 -208 220 -207
rect 220 -208 221 -207
rect 221 -208 222 -207
rect 222 -208 223 -207
rect 223 -208 224 -207
rect 224 -208 225 -207
rect 225 -208 226 -207
rect 226 -208 227 -207
rect 227 -208 228 -207
rect 228 -208 229 -207
rect 229 -208 230 -207
rect 230 -208 231 -207
rect 231 -208 232 -207
rect 232 -208 233 -207
rect 233 -208 234 -207
rect 234 -208 235 -207
rect 235 -208 236 -207
rect 236 -208 237 -207
rect 237 -208 238 -207
rect 238 -208 239 -207
rect 239 -208 240 -207
rect 240 -208 241 -207
rect 241 -208 242 -207
rect 242 -208 243 -207
rect 243 -208 244 -207
rect 244 -208 245 -207
rect 245 -208 246 -207
rect 246 -208 247 -207
rect 247 -208 248 -207
rect 248 -208 249 -207
rect 249 -208 250 -207
rect 250 -208 251 -207
rect 251 -208 252 -207
rect 252 -208 253 -207
rect 253 -208 254 -207
rect 254 -208 255 -207
rect 255 -208 256 -207
rect 256 -208 257 -207
rect 257 -208 258 -207
rect 258 -208 259 -207
rect 259 -208 260 -207
rect 260 -208 261 -207
rect 261 -208 262 -207
rect 262 -208 263 -207
rect 263 -208 264 -207
rect 264 -208 265 -207
rect 265 -208 266 -207
rect 266 -208 267 -207
rect 267 -208 268 -207
rect 268 -208 269 -207
rect 269 -208 270 -207
rect 270 -208 271 -207
rect 271 -208 272 -207
rect 272 -208 273 -207
rect 273 -208 274 -207
rect 274 -208 275 -207
rect 275 -208 276 -207
rect 276 -208 277 -207
rect 277 -208 278 -207
rect 278 -208 279 -207
rect 279 -208 280 -207
rect 280 -208 281 -207
rect 281 -208 282 -207
rect 282 -208 283 -207
rect 283 -208 284 -207
rect 284 -208 285 -207
rect 285 -208 286 -207
rect 286 -208 287 -207
rect 287 -208 288 -207
rect 288 -208 289 -207
rect 289 -208 290 -207
rect 290 -208 291 -207
rect 291 -208 292 -207
rect 292 -208 293 -207
rect 293 -208 294 -207
rect 294 -208 295 -207
rect 295 -208 296 -207
rect 296 -208 297 -207
rect 297 -208 298 -207
rect 298 -208 299 -207
rect 299 -208 300 -207
rect 300 -208 301 -207
rect 301 -208 302 -207
rect 302 -208 303 -207
rect 303 -208 304 -207
rect 304 -208 305 -207
rect 305 -208 306 -207
rect 306 -208 307 -207
rect 307 -208 308 -207
rect 308 -208 309 -207
rect 309 -208 310 -207
rect 310 -208 311 -207
rect 311 -208 312 -207
rect 312 -208 313 -207
rect 313 -208 314 -207
rect 314 -208 315 -207
rect 315 -208 316 -207
rect 316 -208 317 -207
rect 317 -208 318 -207
rect 318 -208 319 -207
rect 319 -208 320 -207
rect 320 -208 321 -207
rect 321 -208 322 -207
rect 322 -208 323 -207
rect 323 -208 324 -207
rect 324 -208 325 -207
rect 325 -208 326 -207
rect 326 -208 327 -207
rect 327 -208 328 -207
rect 328 -208 329 -207
rect 329 -208 330 -207
rect 330 -208 331 -207
rect 331 -208 332 -207
rect 332 -208 333 -207
rect 333 -208 334 -207
rect 334 -208 335 -207
rect 335 -208 336 -207
rect 336 -208 337 -207
rect 337 -208 338 -207
rect 338 -208 339 -207
rect 339 -208 340 -207
rect 340 -208 341 -207
rect 341 -208 342 -207
rect 342 -208 343 -207
rect 343 -208 344 -207
rect 344 -208 345 -207
rect 345 -208 346 -207
rect 346 -208 347 -207
rect 347 -208 348 -207
rect 348 -208 349 -207
rect 349 -208 350 -207
rect 350 -208 351 -207
rect 351 -208 352 -207
rect 352 -208 353 -207
rect 353 -208 354 -207
rect 354 -208 355 -207
rect 355 -208 356 -207
rect 356 -208 357 -207
rect 357 -208 358 -207
rect 358 -208 359 -207
rect 359 -208 360 -207
rect 360 -208 361 -207
rect 361 -208 362 -207
rect 362 -208 363 -207
rect 363 -208 364 -207
rect 364 -208 365 -207
rect 365 -208 366 -207
rect 366 -208 367 -207
rect 367 -208 368 -207
rect 368 -208 369 -207
rect 369 -208 370 -207
rect 370 -208 371 -207
rect 371 -208 372 -207
rect 372 -208 373 -207
rect 373 -208 374 -207
rect 374 -208 375 -207
rect 375 -208 376 -207
rect 376 -208 377 -207
rect 377 -208 378 -207
rect 378 -208 379 -207
rect 379 -208 380 -207
rect 380 -208 381 -207
rect 381 -208 382 -207
rect 382 -208 383 -207
rect 383 -208 384 -207
rect 384 -208 385 -207
rect 385 -208 386 -207
rect 386 -208 387 -207
rect 387 -208 388 -207
rect 388 -208 389 -207
rect 389 -208 390 -207
rect 390 -208 391 -207
rect 391 -208 392 -207
rect 392 -208 393 -207
rect 393 -208 394 -207
rect 394 -208 395 -207
rect 395 -208 396 -207
rect 396 -208 397 -207
rect 397 -208 398 -207
rect 398 -208 399 -207
rect 399 -208 400 -207
rect 400 -208 401 -207
rect 401 -208 402 -207
rect 402 -208 403 -207
rect 403 -208 404 -207
rect 404 -208 405 -207
rect 405 -208 406 -207
rect 406 -208 407 -207
rect 407 -208 408 -207
rect 408 -208 409 -207
rect 409 -208 410 -207
rect 410 -208 411 -207
rect 411 -208 412 -207
rect 412 -208 413 -207
rect 413 -208 414 -207
rect 414 -208 415 -207
rect 415 -208 416 -207
rect 416 -208 417 -207
rect 417 -208 418 -207
rect 418 -208 419 -207
rect 419 -208 420 -207
rect 420 -208 421 -207
rect 421 -208 422 -207
rect 422 -208 423 -207
rect 423 -208 424 -207
rect 424 -208 425 -207
rect 425 -208 426 -207
rect 426 -208 427 -207
rect 427 -208 428 -207
rect 428 -208 429 -207
rect 429 -208 430 -207
rect 430 -208 431 -207
rect 431 -208 432 -207
rect 432 -208 433 -207
rect 433 -208 434 -207
rect 434 -208 435 -207
rect 435 -208 436 -207
rect 436 -208 437 -207
rect 437 -208 438 -207
rect 438 -208 439 -207
rect 439 -208 440 -207
rect 440 -208 441 -207
rect 441 -208 442 -207
rect 442 -208 443 -207
rect 443 -208 444 -207
rect 444 -208 445 -207
rect 445 -208 446 -207
rect 446 -208 447 -207
rect 447 -208 448 -207
rect 448 -208 449 -207
rect 449 -208 450 -207
rect 450 -208 451 -207
rect 451 -208 452 -207
rect 452 -208 453 -207
rect 453 -208 454 -207
rect 454 -208 455 -207
rect 455 -208 456 -207
rect 456 -208 457 -207
rect 457 -208 458 -207
rect 458 -208 459 -207
rect 459 -208 460 -207
rect 460 -208 461 -207
rect 461 -208 462 -207
rect 462 -208 463 -207
rect 463 -208 464 -207
rect 464 -208 465 -207
rect 465 -208 466 -207
rect 466 -208 467 -207
rect 467 -208 468 -207
rect 468 -208 469 -207
rect 469 -208 470 -207
rect 470 -208 471 -207
rect 471 -208 472 -207
rect 472 -208 473 -207
rect 473 -208 474 -207
rect 474 -208 475 -207
rect 475 -208 476 -207
rect 476 -208 477 -207
rect 477 -208 478 -207
rect 478 -208 479 -207
rect 479 -208 480 -207
rect 2 -209 3 -208
rect 3 -209 4 -208
rect 4 -209 5 -208
rect 5 -209 6 -208
rect 6 -209 7 -208
rect 7 -209 8 -208
rect 8 -209 9 -208
rect 9 -209 10 -208
rect 10 -209 11 -208
rect 11 -209 12 -208
rect 12 -209 13 -208
rect 13 -209 14 -208
rect 14 -209 15 -208
rect 15 -209 16 -208
rect 16 -209 17 -208
rect 17 -209 18 -208
rect 18 -209 19 -208
rect 19 -209 20 -208
rect 20 -209 21 -208
rect 21 -209 22 -208
rect 22 -209 23 -208
rect 23 -209 24 -208
rect 24 -209 25 -208
rect 25 -209 26 -208
rect 26 -209 27 -208
rect 27 -209 28 -208
rect 28 -209 29 -208
rect 29 -209 30 -208
rect 30 -209 31 -208
rect 31 -209 32 -208
rect 32 -209 33 -208
rect 33 -209 34 -208
rect 34 -209 35 -208
rect 35 -209 36 -208
rect 36 -209 37 -208
rect 37 -209 38 -208
rect 38 -209 39 -208
rect 39 -209 40 -208
rect 40 -209 41 -208
rect 41 -209 42 -208
rect 42 -209 43 -208
rect 43 -209 44 -208
rect 44 -209 45 -208
rect 45 -209 46 -208
rect 46 -209 47 -208
rect 47 -209 48 -208
rect 48 -209 49 -208
rect 49 -209 50 -208
rect 50 -209 51 -208
rect 51 -209 52 -208
rect 52 -209 53 -208
rect 53 -209 54 -208
rect 54 -209 55 -208
rect 55 -209 56 -208
rect 56 -209 57 -208
rect 57 -209 58 -208
rect 58 -209 59 -208
rect 59 -209 60 -208
rect 60 -209 61 -208
rect 61 -209 62 -208
rect 62 -209 63 -208
rect 63 -209 64 -208
rect 64 -209 65 -208
rect 65 -209 66 -208
rect 66 -209 67 -208
rect 67 -209 68 -208
rect 68 -209 69 -208
rect 69 -209 70 -208
rect 70 -209 71 -208
rect 71 -209 72 -208
rect 72 -209 73 -208
rect 73 -209 74 -208
rect 74 -209 75 -208
rect 75 -209 76 -208
rect 76 -209 77 -208
rect 77 -209 78 -208
rect 78 -209 79 -208
rect 79 -209 80 -208
rect 80 -209 81 -208
rect 81 -209 82 -208
rect 82 -209 83 -208
rect 83 -209 84 -208
rect 84 -209 85 -208
rect 85 -209 86 -208
rect 86 -209 87 -208
rect 87 -209 88 -208
rect 88 -209 89 -208
rect 89 -209 90 -208
rect 90 -209 91 -208
rect 91 -209 92 -208
rect 92 -209 93 -208
rect 93 -209 94 -208
rect 94 -209 95 -208
rect 95 -209 96 -208
rect 96 -209 97 -208
rect 97 -209 98 -208
rect 98 -209 99 -208
rect 99 -209 100 -208
rect 100 -209 101 -208
rect 101 -209 102 -208
rect 102 -209 103 -208
rect 103 -209 104 -208
rect 104 -209 105 -208
rect 105 -209 106 -208
rect 106 -209 107 -208
rect 107 -209 108 -208
rect 108 -209 109 -208
rect 109 -209 110 -208
rect 110 -209 111 -208
rect 111 -209 112 -208
rect 112 -209 113 -208
rect 113 -209 114 -208
rect 114 -209 115 -208
rect 115 -209 116 -208
rect 116 -209 117 -208
rect 117 -209 118 -208
rect 118 -209 119 -208
rect 119 -209 120 -208
rect 120 -209 121 -208
rect 121 -209 122 -208
rect 122 -209 123 -208
rect 123 -209 124 -208
rect 124 -209 125 -208
rect 125 -209 126 -208
rect 126 -209 127 -208
rect 127 -209 128 -208
rect 128 -209 129 -208
rect 129 -209 130 -208
rect 130 -209 131 -208
rect 131 -209 132 -208
rect 132 -209 133 -208
rect 133 -209 134 -208
rect 134 -209 135 -208
rect 135 -209 136 -208
rect 136 -209 137 -208
rect 137 -209 138 -208
rect 138 -209 139 -208
rect 139 -209 140 -208
rect 140 -209 141 -208
rect 141 -209 142 -208
rect 142 -209 143 -208
rect 143 -209 144 -208
rect 144 -209 145 -208
rect 145 -209 146 -208
rect 146 -209 147 -208
rect 147 -209 148 -208
rect 148 -209 149 -208
rect 149 -209 150 -208
rect 150 -209 151 -208
rect 151 -209 152 -208
rect 152 -209 153 -208
rect 153 -209 154 -208
rect 154 -209 155 -208
rect 155 -209 156 -208
rect 156 -209 157 -208
rect 157 -209 158 -208
rect 158 -209 159 -208
rect 159 -209 160 -208
rect 160 -209 161 -208
rect 161 -209 162 -208
rect 162 -209 163 -208
rect 163 -209 164 -208
rect 164 -209 165 -208
rect 165 -209 166 -208
rect 166 -209 167 -208
rect 167 -209 168 -208
rect 168 -209 169 -208
rect 169 -209 170 -208
rect 170 -209 171 -208
rect 171 -209 172 -208
rect 172 -209 173 -208
rect 173 -209 174 -208
rect 174 -209 175 -208
rect 175 -209 176 -208
rect 176 -209 177 -208
rect 177 -209 178 -208
rect 178 -209 179 -208
rect 179 -209 180 -208
rect 180 -209 181 -208
rect 181 -209 182 -208
rect 182 -209 183 -208
rect 183 -209 184 -208
rect 184 -209 185 -208
rect 185 -209 186 -208
rect 186 -209 187 -208
rect 187 -209 188 -208
rect 188 -209 189 -208
rect 189 -209 190 -208
rect 190 -209 191 -208
rect 191 -209 192 -208
rect 192 -209 193 -208
rect 193 -209 194 -208
rect 194 -209 195 -208
rect 195 -209 196 -208
rect 196 -209 197 -208
rect 197 -209 198 -208
rect 198 -209 199 -208
rect 199 -209 200 -208
rect 200 -209 201 -208
rect 201 -209 202 -208
rect 202 -209 203 -208
rect 203 -209 204 -208
rect 204 -209 205 -208
rect 205 -209 206 -208
rect 206 -209 207 -208
rect 207 -209 208 -208
rect 208 -209 209 -208
rect 209 -209 210 -208
rect 210 -209 211 -208
rect 211 -209 212 -208
rect 212 -209 213 -208
rect 213 -209 214 -208
rect 214 -209 215 -208
rect 215 -209 216 -208
rect 216 -209 217 -208
rect 217 -209 218 -208
rect 218 -209 219 -208
rect 219 -209 220 -208
rect 220 -209 221 -208
rect 221 -209 222 -208
rect 222 -209 223 -208
rect 223 -209 224 -208
rect 224 -209 225 -208
rect 225 -209 226 -208
rect 226 -209 227 -208
rect 227 -209 228 -208
rect 228 -209 229 -208
rect 229 -209 230 -208
rect 230 -209 231 -208
rect 231 -209 232 -208
rect 232 -209 233 -208
rect 233 -209 234 -208
rect 234 -209 235 -208
rect 235 -209 236 -208
rect 236 -209 237 -208
rect 237 -209 238 -208
rect 238 -209 239 -208
rect 239 -209 240 -208
rect 240 -209 241 -208
rect 241 -209 242 -208
rect 242 -209 243 -208
rect 243 -209 244 -208
rect 244 -209 245 -208
rect 245 -209 246 -208
rect 246 -209 247 -208
rect 247 -209 248 -208
rect 248 -209 249 -208
rect 249 -209 250 -208
rect 250 -209 251 -208
rect 251 -209 252 -208
rect 252 -209 253 -208
rect 253 -209 254 -208
rect 254 -209 255 -208
rect 255 -209 256 -208
rect 256 -209 257 -208
rect 257 -209 258 -208
rect 258 -209 259 -208
rect 259 -209 260 -208
rect 260 -209 261 -208
rect 261 -209 262 -208
rect 262 -209 263 -208
rect 263 -209 264 -208
rect 264 -209 265 -208
rect 265 -209 266 -208
rect 266 -209 267 -208
rect 267 -209 268 -208
rect 268 -209 269 -208
rect 269 -209 270 -208
rect 270 -209 271 -208
rect 271 -209 272 -208
rect 272 -209 273 -208
rect 273 -209 274 -208
rect 274 -209 275 -208
rect 275 -209 276 -208
rect 276 -209 277 -208
rect 277 -209 278 -208
rect 278 -209 279 -208
rect 279 -209 280 -208
rect 280 -209 281 -208
rect 281 -209 282 -208
rect 282 -209 283 -208
rect 283 -209 284 -208
rect 284 -209 285 -208
rect 285 -209 286 -208
rect 286 -209 287 -208
rect 287 -209 288 -208
rect 288 -209 289 -208
rect 289 -209 290 -208
rect 290 -209 291 -208
rect 291 -209 292 -208
rect 292 -209 293 -208
rect 293 -209 294 -208
rect 294 -209 295 -208
rect 295 -209 296 -208
rect 296 -209 297 -208
rect 297 -209 298 -208
rect 298 -209 299 -208
rect 299 -209 300 -208
rect 300 -209 301 -208
rect 301 -209 302 -208
rect 302 -209 303 -208
rect 303 -209 304 -208
rect 304 -209 305 -208
rect 305 -209 306 -208
rect 306 -209 307 -208
rect 307 -209 308 -208
rect 308 -209 309 -208
rect 309 -209 310 -208
rect 310 -209 311 -208
rect 311 -209 312 -208
rect 312 -209 313 -208
rect 313 -209 314 -208
rect 314 -209 315 -208
rect 315 -209 316 -208
rect 316 -209 317 -208
rect 317 -209 318 -208
rect 318 -209 319 -208
rect 319 -209 320 -208
rect 320 -209 321 -208
rect 321 -209 322 -208
rect 322 -209 323 -208
rect 323 -209 324 -208
rect 324 -209 325 -208
rect 325 -209 326 -208
rect 326 -209 327 -208
rect 327 -209 328 -208
rect 328 -209 329 -208
rect 329 -209 330 -208
rect 330 -209 331 -208
rect 331 -209 332 -208
rect 332 -209 333 -208
rect 333 -209 334 -208
rect 334 -209 335 -208
rect 335 -209 336 -208
rect 336 -209 337 -208
rect 337 -209 338 -208
rect 338 -209 339 -208
rect 339 -209 340 -208
rect 340 -209 341 -208
rect 341 -209 342 -208
rect 342 -209 343 -208
rect 343 -209 344 -208
rect 344 -209 345 -208
rect 345 -209 346 -208
rect 346 -209 347 -208
rect 347 -209 348 -208
rect 348 -209 349 -208
rect 349 -209 350 -208
rect 350 -209 351 -208
rect 351 -209 352 -208
rect 352 -209 353 -208
rect 353 -209 354 -208
rect 354 -209 355 -208
rect 355 -209 356 -208
rect 356 -209 357 -208
rect 357 -209 358 -208
rect 358 -209 359 -208
rect 359 -209 360 -208
rect 360 -209 361 -208
rect 361 -209 362 -208
rect 362 -209 363 -208
rect 363 -209 364 -208
rect 364 -209 365 -208
rect 365 -209 366 -208
rect 366 -209 367 -208
rect 367 -209 368 -208
rect 368 -209 369 -208
rect 369 -209 370 -208
rect 370 -209 371 -208
rect 371 -209 372 -208
rect 372 -209 373 -208
rect 373 -209 374 -208
rect 374 -209 375 -208
rect 375 -209 376 -208
rect 376 -209 377 -208
rect 377 -209 378 -208
rect 378 -209 379 -208
rect 379 -209 380 -208
rect 380 -209 381 -208
rect 381 -209 382 -208
rect 382 -209 383 -208
rect 383 -209 384 -208
rect 384 -209 385 -208
rect 385 -209 386 -208
rect 386 -209 387 -208
rect 387 -209 388 -208
rect 388 -209 389 -208
rect 389 -209 390 -208
rect 390 -209 391 -208
rect 391 -209 392 -208
rect 392 -209 393 -208
rect 393 -209 394 -208
rect 394 -209 395 -208
rect 395 -209 396 -208
rect 396 -209 397 -208
rect 397 -209 398 -208
rect 398 -209 399 -208
rect 399 -209 400 -208
rect 400 -209 401 -208
rect 401 -209 402 -208
rect 402 -209 403 -208
rect 403 -209 404 -208
rect 404 -209 405 -208
rect 405 -209 406 -208
rect 406 -209 407 -208
rect 407 -209 408 -208
rect 408 -209 409 -208
rect 409 -209 410 -208
rect 410 -209 411 -208
rect 411 -209 412 -208
rect 412 -209 413 -208
rect 413 -209 414 -208
rect 414 -209 415 -208
rect 415 -209 416 -208
rect 416 -209 417 -208
rect 417 -209 418 -208
rect 418 -209 419 -208
rect 419 -209 420 -208
rect 420 -209 421 -208
rect 421 -209 422 -208
rect 422 -209 423 -208
rect 423 -209 424 -208
rect 424 -209 425 -208
rect 425 -209 426 -208
rect 426 -209 427 -208
rect 427 -209 428 -208
rect 428 -209 429 -208
rect 429 -209 430 -208
rect 430 -209 431 -208
rect 431 -209 432 -208
rect 432 -209 433 -208
rect 433 -209 434 -208
rect 434 -209 435 -208
rect 435 -209 436 -208
rect 436 -209 437 -208
rect 437 -209 438 -208
rect 438 -209 439 -208
rect 439 -209 440 -208
rect 440 -209 441 -208
rect 441 -209 442 -208
rect 442 -209 443 -208
rect 443 -209 444 -208
rect 444 -209 445 -208
rect 445 -209 446 -208
rect 446 -209 447 -208
rect 447 -209 448 -208
rect 448 -209 449 -208
rect 449 -209 450 -208
rect 450 -209 451 -208
rect 451 -209 452 -208
rect 452 -209 453 -208
rect 453 -209 454 -208
rect 454 -209 455 -208
rect 455 -209 456 -208
rect 456 -209 457 -208
rect 457 -209 458 -208
rect 458 -209 459 -208
rect 459 -209 460 -208
rect 460 -209 461 -208
rect 461 -209 462 -208
rect 462 -209 463 -208
rect 463 -209 464 -208
rect 464 -209 465 -208
rect 465 -209 466 -208
rect 466 -209 467 -208
rect 467 -209 468 -208
rect 468 -209 469 -208
rect 469 -209 470 -208
rect 470 -209 471 -208
rect 471 -209 472 -208
rect 472 -209 473 -208
rect 473 -209 474 -208
rect 474 -209 475 -208
rect 475 -209 476 -208
rect 476 -209 477 -208
rect 477 -209 478 -208
rect 478 -209 479 -208
rect 479 -209 480 -208
rect 2 -210 3 -209
rect 3 -210 4 -209
rect 4 -210 5 -209
rect 5 -210 6 -209
rect 6 -210 7 -209
rect 7 -210 8 -209
rect 8 -210 9 -209
rect 9 -210 10 -209
rect 10 -210 11 -209
rect 11 -210 12 -209
rect 12 -210 13 -209
rect 13 -210 14 -209
rect 14 -210 15 -209
rect 15 -210 16 -209
rect 16 -210 17 -209
rect 17 -210 18 -209
rect 18 -210 19 -209
rect 19 -210 20 -209
rect 20 -210 21 -209
rect 21 -210 22 -209
rect 22 -210 23 -209
rect 23 -210 24 -209
rect 24 -210 25 -209
rect 25 -210 26 -209
rect 26 -210 27 -209
rect 27 -210 28 -209
rect 28 -210 29 -209
rect 29 -210 30 -209
rect 30 -210 31 -209
rect 31 -210 32 -209
rect 32 -210 33 -209
rect 33 -210 34 -209
rect 34 -210 35 -209
rect 35 -210 36 -209
rect 36 -210 37 -209
rect 37 -210 38 -209
rect 38 -210 39 -209
rect 39 -210 40 -209
rect 40 -210 41 -209
rect 41 -210 42 -209
rect 42 -210 43 -209
rect 43 -210 44 -209
rect 44 -210 45 -209
rect 45 -210 46 -209
rect 46 -210 47 -209
rect 47 -210 48 -209
rect 48 -210 49 -209
rect 49 -210 50 -209
rect 50 -210 51 -209
rect 51 -210 52 -209
rect 52 -210 53 -209
rect 53 -210 54 -209
rect 54 -210 55 -209
rect 55 -210 56 -209
rect 56 -210 57 -209
rect 57 -210 58 -209
rect 58 -210 59 -209
rect 59 -210 60 -209
rect 60 -210 61 -209
rect 61 -210 62 -209
rect 62 -210 63 -209
rect 63 -210 64 -209
rect 64 -210 65 -209
rect 65 -210 66 -209
rect 66 -210 67 -209
rect 67 -210 68 -209
rect 68 -210 69 -209
rect 69 -210 70 -209
rect 70 -210 71 -209
rect 71 -210 72 -209
rect 72 -210 73 -209
rect 73 -210 74 -209
rect 74 -210 75 -209
rect 75 -210 76 -209
rect 76 -210 77 -209
rect 77 -210 78 -209
rect 78 -210 79 -209
rect 79 -210 80 -209
rect 80 -210 81 -209
rect 81 -210 82 -209
rect 82 -210 83 -209
rect 83 -210 84 -209
rect 84 -210 85 -209
rect 85 -210 86 -209
rect 86 -210 87 -209
rect 87 -210 88 -209
rect 88 -210 89 -209
rect 89 -210 90 -209
rect 90 -210 91 -209
rect 91 -210 92 -209
rect 92 -210 93 -209
rect 93 -210 94 -209
rect 94 -210 95 -209
rect 95 -210 96 -209
rect 96 -210 97 -209
rect 97 -210 98 -209
rect 98 -210 99 -209
rect 99 -210 100 -209
rect 100 -210 101 -209
rect 101 -210 102 -209
rect 102 -210 103 -209
rect 103 -210 104 -209
rect 104 -210 105 -209
rect 105 -210 106 -209
rect 106 -210 107 -209
rect 107 -210 108 -209
rect 108 -210 109 -209
rect 109 -210 110 -209
rect 110 -210 111 -209
rect 111 -210 112 -209
rect 112 -210 113 -209
rect 113 -210 114 -209
rect 114 -210 115 -209
rect 115 -210 116 -209
rect 116 -210 117 -209
rect 117 -210 118 -209
rect 118 -210 119 -209
rect 119 -210 120 -209
rect 120 -210 121 -209
rect 121 -210 122 -209
rect 122 -210 123 -209
rect 123 -210 124 -209
rect 124 -210 125 -209
rect 125 -210 126 -209
rect 126 -210 127 -209
rect 127 -210 128 -209
rect 128 -210 129 -209
rect 129 -210 130 -209
rect 130 -210 131 -209
rect 131 -210 132 -209
rect 132 -210 133 -209
rect 133 -210 134 -209
rect 134 -210 135 -209
rect 135 -210 136 -209
rect 136 -210 137 -209
rect 137 -210 138 -209
rect 138 -210 139 -209
rect 139 -210 140 -209
rect 140 -210 141 -209
rect 141 -210 142 -209
rect 142 -210 143 -209
rect 143 -210 144 -209
rect 144 -210 145 -209
rect 145 -210 146 -209
rect 146 -210 147 -209
rect 147 -210 148 -209
rect 148 -210 149 -209
rect 149 -210 150 -209
rect 150 -210 151 -209
rect 151 -210 152 -209
rect 152 -210 153 -209
rect 153 -210 154 -209
rect 154 -210 155 -209
rect 155 -210 156 -209
rect 156 -210 157 -209
rect 157 -210 158 -209
rect 158 -210 159 -209
rect 159 -210 160 -209
rect 160 -210 161 -209
rect 161 -210 162 -209
rect 162 -210 163 -209
rect 163 -210 164 -209
rect 164 -210 165 -209
rect 165 -210 166 -209
rect 166 -210 167 -209
rect 167 -210 168 -209
rect 168 -210 169 -209
rect 169 -210 170 -209
rect 170 -210 171 -209
rect 171 -210 172 -209
rect 172 -210 173 -209
rect 173 -210 174 -209
rect 174 -210 175 -209
rect 175 -210 176 -209
rect 176 -210 177 -209
rect 177 -210 178 -209
rect 178 -210 179 -209
rect 179 -210 180 -209
rect 180 -210 181 -209
rect 181 -210 182 -209
rect 182 -210 183 -209
rect 183 -210 184 -209
rect 184 -210 185 -209
rect 185 -210 186 -209
rect 186 -210 187 -209
rect 187 -210 188 -209
rect 188 -210 189 -209
rect 189 -210 190 -209
rect 190 -210 191 -209
rect 191 -210 192 -209
rect 192 -210 193 -209
rect 193 -210 194 -209
rect 194 -210 195 -209
rect 195 -210 196 -209
rect 196 -210 197 -209
rect 197 -210 198 -209
rect 198 -210 199 -209
rect 199 -210 200 -209
rect 200 -210 201 -209
rect 201 -210 202 -209
rect 202 -210 203 -209
rect 203 -210 204 -209
rect 204 -210 205 -209
rect 205 -210 206 -209
rect 206 -210 207 -209
rect 207 -210 208 -209
rect 208 -210 209 -209
rect 209 -210 210 -209
rect 210 -210 211 -209
rect 211 -210 212 -209
rect 212 -210 213 -209
rect 213 -210 214 -209
rect 214 -210 215 -209
rect 215 -210 216 -209
rect 216 -210 217 -209
rect 217 -210 218 -209
rect 218 -210 219 -209
rect 219 -210 220 -209
rect 220 -210 221 -209
rect 221 -210 222 -209
rect 222 -210 223 -209
rect 223 -210 224 -209
rect 224 -210 225 -209
rect 225 -210 226 -209
rect 226 -210 227 -209
rect 227 -210 228 -209
rect 228 -210 229 -209
rect 229 -210 230 -209
rect 230 -210 231 -209
rect 231 -210 232 -209
rect 232 -210 233 -209
rect 233 -210 234 -209
rect 234 -210 235 -209
rect 235 -210 236 -209
rect 236 -210 237 -209
rect 237 -210 238 -209
rect 238 -210 239 -209
rect 239 -210 240 -209
rect 240 -210 241 -209
rect 241 -210 242 -209
rect 242 -210 243 -209
rect 243 -210 244 -209
rect 244 -210 245 -209
rect 245 -210 246 -209
rect 246 -210 247 -209
rect 247 -210 248 -209
rect 248 -210 249 -209
rect 249 -210 250 -209
rect 250 -210 251 -209
rect 251 -210 252 -209
rect 252 -210 253 -209
rect 253 -210 254 -209
rect 254 -210 255 -209
rect 255 -210 256 -209
rect 256 -210 257 -209
rect 257 -210 258 -209
rect 258 -210 259 -209
rect 259 -210 260 -209
rect 260 -210 261 -209
rect 261 -210 262 -209
rect 262 -210 263 -209
rect 263 -210 264 -209
rect 264 -210 265 -209
rect 265 -210 266 -209
rect 266 -210 267 -209
rect 267 -210 268 -209
rect 268 -210 269 -209
rect 269 -210 270 -209
rect 270 -210 271 -209
rect 271 -210 272 -209
rect 272 -210 273 -209
rect 273 -210 274 -209
rect 274 -210 275 -209
rect 275 -210 276 -209
rect 276 -210 277 -209
rect 277 -210 278 -209
rect 278 -210 279 -209
rect 279 -210 280 -209
rect 280 -210 281 -209
rect 281 -210 282 -209
rect 282 -210 283 -209
rect 283 -210 284 -209
rect 284 -210 285 -209
rect 285 -210 286 -209
rect 286 -210 287 -209
rect 287 -210 288 -209
rect 288 -210 289 -209
rect 289 -210 290 -209
rect 290 -210 291 -209
rect 291 -210 292 -209
rect 292 -210 293 -209
rect 293 -210 294 -209
rect 294 -210 295 -209
rect 295 -210 296 -209
rect 296 -210 297 -209
rect 297 -210 298 -209
rect 298 -210 299 -209
rect 299 -210 300 -209
rect 300 -210 301 -209
rect 301 -210 302 -209
rect 302 -210 303 -209
rect 303 -210 304 -209
rect 304 -210 305 -209
rect 305 -210 306 -209
rect 306 -210 307 -209
rect 307 -210 308 -209
rect 308 -210 309 -209
rect 309 -210 310 -209
rect 310 -210 311 -209
rect 311 -210 312 -209
rect 312 -210 313 -209
rect 313 -210 314 -209
rect 314 -210 315 -209
rect 315 -210 316 -209
rect 316 -210 317 -209
rect 317 -210 318 -209
rect 318 -210 319 -209
rect 319 -210 320 -209
rect 320 -210 321 -209
rect 321 -210 322 -209
rect 322 -210 323 -209
rect 323 -210 324 -209
rect 324 -210 325 -209
rect 325 -210 326 -209
rect 326 -210 327 -209
rect 327 -210 328 -209
rect 328 -210 329 -209
rect 329 -210 330 -209
rect 330 -210 331 -209
rect 331 -210 332 -209
rect 332 -210 333 -209
rect 333 -210 334 -209
rect 334 -210 335 -209
rect 335 -210 336 -209
rect 336 -210 337 -209
rect 337 -210 338 -209
rect 338 -210 339 -209
rect 339 -210 340 -209
rect 340 -210 341 -209
rect 341 -210 342 -209
rect 342 -210 343 -209
rect 343 -210 344 -209
rect 344 -210 345 -209
rect 345 -210 346 -209
rect 346 -210 347 -209
rect 347 -210 348 -209
rect 348 -210 349 -209
rect 349 -210 350 -209
rect 350 -210 351 -209
rect 351 -210 352 -209
rect 352 -210 353 -209
rect 353 -210 354 -209
rect 354 -210 355 -209
rect 355 -210 356 -209
rect 356 -210 357 -209
rect 357 -210 358 -209
rect 358 -210 359 -209
rect 359 -210 360 -209
rect 360 -210 361 -209
rect 361 -210 362 -209
rect 362 -210 363 -209
rect 363 -210 364 -209
rect 364 -210 365 -209
rect 365 -210 366 -209
rect 366 -210 367 -209
rect 367 -210 368 -209
rect 368 -210 369 -209
rect 369 -210 370 -209
rect 370 -210 371 -209
rect 371 -210 372 -209
rect 372 -210 373 -209
rect 373 -210 374 -209
rect 374 -210 375 -209
rect 375 -210 376 -209
rect 376 -210 377 -209
rect 377 -210 378 -209
rect 378 -210 379 -209
rect 379 -210 380 -209
rect 380 -210 381 -209
rect 381 -210 382 -209
rect 382 -210 383 -209
rect 383 -210 384 -209
rect 384 -210 385 -209
rect 385 -210 386 -209
rect 386 -210 387 -209
rect 387 -210 388 -209
rect 388 -210 389 -209
rect 389 -210 390 -209
rect 390 -210 391 -209
rect 391 -210 392 -209
rect 392 -210 393 -209
rect 393 -210 394 -209
rect 394 -210 395 -209
rect 395 -210 396 -209
rect 396 -210 397 -209
rect 397 -210 398 -209
rect 398 -210 399 -209
rect 399 -210 400 -209
rect 400 -210 401 -209
rect 401 -210 402 -209
rect 402 -210 403 -209
rect 403 -210 404 -209
rect 404 -210 405 -209
rect 405 -210 406 -209
rect 406 -210 407 -209
rect 407 -210 408 -209
rect 408 -210 409 -209
rect 409 -210 410 -209
rect 410 -210 411 -209
rect 411 -210 412 -209
rect 412 -210 413 -209
rect 413 -210 414 -209
rect 414 -210 415 -209
rect 415 -210 416 -209
rect 416 -210 417 -209
rect 417 -210 418 -209
rect 418 -210 419 -209
rect 419 -210 420 -209
rect 420 -210 421 -209
rect 421 -210 422 -209
rect 422 -210 423 -209
rect 423 -210 424 -209
rect 424 -210 425 -209
rect 425 -210 426 -209
rect 426 -210 427 -209
rect 427 -210 428 -209
rect 428 -210 429 -209
rect 429 -210 430 -209
rect 430 -210 431 -209
rect 431 -210 432 -209
rect 432 -210 433 -209
rect 433 -210 434 -209
rect 434 -210 435 -209
rect 435 -210 436 -209
rect 436 -210 437 -209
rect 437 -210 438 -209
rect 438 -210 439 -209
rect 439 -210 440 -209
rect 440 -210 441 -209
rect 441 -210 442 -209
rect 442 -210 443 -209
rect 443 -210 444 -209
rect 444 -210 445 -209
rect 445 -210 446 -209
rect 446 -210 447 -209
rect 447 -210 448 -209
rect 448 -210 449 -209
rect 449 -210 450 -209
rect 450 -210 451 -209
rect 451 -210 452 -209
rect 452 -210 453 -209
rect 453 -210 454 -209
rect 454 -210 455 -209
rect 455 -210 456 -209
rect 456 -210 457 -209
rect 457 -210 458 -209
rect 458 -210 459 -209
rect 459 -210 460 -209
rect 460 -210 461 -209
rect 461 -210 462 -209
rect 462 -210 463 -209
rect 463 -210 464 -209
rect 464 -210 465 -209
rect 465 -210 466 -209
rect 466 -210 467 -209
rect 467 -210 468 -209
rect 468 -210 469 -209
rect 469 -210 470 -209
rect 470 -210 471 -209
rect 471 -210 472 -209
rect 472 -210 473 -209
rect 473 -210 474 -209
rect 474 -210 475 -209
rect 475 -210 476 -209
rect 476 -210 477 -209
rect 477 -210 478 -209
rect 478 -210 479 -209
rect 479 -210 480 -209
rect 2 -211 3 -210
rect 3 -211 4 -210
rect 4 -211 5 -210
rect 5 -211 6 -210
rect 6 -211 7 -210
rect 7 -211 8 -210
rect 8 -211 9 -210
rect 9 -211 10 -210
rect 10 -211 11 -210
rect 11 -211 12 -210
rect 12 -211 13 -210
rect 13 -211 14 -210
rect 14 -211 15 -210
rect 15 -211 16 -210
rect 16 -211 17 -210
rect 17 -211 18 -210
rect 18 -211 19 -210
rect 19 -211 20 -210
rect 20 -211 21 -210
rect 21 -211 22 -210
rect 22 -211 23 -210
rect 23 -211 24 -210
rect 24 -211 25 -210
rect 25 -211 26 -210
rect 26 -211 27 -210
rect 27 -211 28 -210
rect 28 -211 29 -210
rect 29 -211 30 -210
rect 30 -211 31 -210
rect 31 -211 32 -210
rect 32 -211 33 -210
rect 33 -211 34 -210
rect 34 -211 35 -210
rect 35 -211 36 -210
rect 36 -211 37 -210
rect 37 -211 38 -210
rect 38 -211 39 -210
rect 39 -211 40 -210
rect 40 -211 41 -210
rect 41 -211 42 -210
rect 42 -211 43 -210
rect 43 -211 44 -210
rect 44 -211 45 -210
rect 45 -211 46 -210
rect 46 -211 47 -210
rect 47 -211 48 -210
rect 48 -211 49 -210
rect 49 -211 50 -210
rect 50 -211 51 -210
rect 51 -211 52 -210
rect 52 -211 53 -210
rect 53 -211 54 -210
rect 54 -211 55 -210
rect 55 -211 56 -210
rect 56 -211 57 -210
rect 57 -211 58 -210
rect 58 -211 59 -210
rect 59 -211 60 -210
rect 60 -211 61 -210
rect 61 -211 62 -210
rect 62 -211 63 -210
rect 63 -211 64 -210
rect 64 -211 65 -210
rect 65 -211 66 -210
rect 66 -211 67 -210
rect 67 -211 68 -210
rect 68 -211 69 -210
rect 69 -211 70 -210
rect 70 -211 71 -210
rect 71 -211 72 -210
rect 72 -211 73 -210
rect 73 -211 74 -210
rect 74 -211 75 -210
rect 75 -211 76 -210
rect 76 -211 77 -210
rect 77 -211 78 -210
rect 78 -211 79 -210
rect 79 -211 80 -210
rect 80 -211 81 -210
rect 81 -211 82 -210
rect 82 -211 83 -210
rect 83 -211 84 -210
rect 84 -211 85 -210
rect 85 -211 86 -210
rect 86 -211 87 -210
rect 87 -211 88 -210
rect 88 -211 89 -210
rect 89 -211 90 -210
rect 90 -211 91 -210
rect 91 -211 92 -210
rect 92 -211 93 -210
rect 93 -211 94 -210
rect 94 -211 95 -210
rect 95 -211 96 -210
rect 96 -211 97 -210
rect 97 -211 98 -210
rect 98 -211 99 -210
rect 99 -211 100 -210
rect 100 -211 101 -210
rect 101 -211 102 -210
rect 102 -211 103 -210
rect 103 -211 104 -210
rect 104 -211 105 -210
rect 105 -211 106 -210
rect 106 -211 107 -210
rect 107 -211 108 -210
rect 108 -211 109 -210
rect 109 -211 110 -210
rect 110 -211 111 -210
rect 111 -211 112 -210
rect 112 -211 113 -210
rect 113 -211 114 -210
rect 114 -211 115 -210
rect 115 -211 116 -210
rect 116 -211 117 -210
rect 117 -211 118 -210
rect 118 -211 119 -210
rect 119 -211 120 -210
rect 120 -211 121 -210
rect 121 -211 122 -210
rect 122 -211 123 -210
rect 123 -211 124 -210
rect 124 -211 125 -210
rect 125 -211 126 -210
rect 126 -211 127 -210
rect 127 -211 128 -210
rect 128 -211 129 -210
rect 129 -211 130 -210
rect 130 -211 131 -210
rect 131 -211 132 -210
rect 132 -211 133 -210
rect 133 -211 134 -210
rect 134 -211 135 -210
rect 135 -211 136 -210
rect 136 -211 137 -210
rect 137 -211 138 -210
rect 138 -211 139 -210
rect 139 -211 140 -210
rect 140 -211 141 -210
rect 141 -211 142 -210
rect 142 -211 143 -210
rect 143 -211 144 -210
rect 144 -211 145 -210
rect 145 -211 146 -210
rect 146 -211 147 -210
rect 147 -211 148 -210
rect 148 -211 149 -210
rect 149 -211 150 -210
rect 150 -211 151 -210
rect 151 -211 152 -210
rect 152 -211 153 -210
rect 153 -211 154 -210
rect 154 -211 155 -210
rect 155 -211 156 -210
rect 156 -211 157 -210
rect 157 -211 158 -210
rect 158 -211 159 -210
rect 159 -211 160 -210
rect 160 -211 161 -210
rect 161 -211 162 -210
rect 162 -211 163 -210
rect 163 -211 164 -210
rect 164 -211 165 -210
rect 165 -211 166 -210
rect 166 -211 167 -210
rect 167 -211 168 -210
rect 168 -211 169 -210
rect 169 -211 170 -210
rect 170 -211 171 -210
rect 171 -211 172 -210
rect 172 -211 173 -210
rect 173 -211 174 -210
rect 174 -211 175 -210
rect 175 -211 176 -210
rect 176 -211 177 -210
rect 177 -211 178 -210
rect 178 -211 179 -210
rect 179 -211 180 -210
rect 180 -211 181 -210
rect 181 -211 182 -210
rect 182 -211 183 -210
rect 183 -211 184 -210
rect 184 -211 185 -210
rect 185 -211 186 -210
rect 186 -211 187 -210
rect 187 -211 188 -210
rect 188 -211 189 -210
rect 189 -211 190 -210
rect 190 -211 191 -210
rect 191 -211 192 -210
rect 192 -211 193 -210
rect 193 -211 194 -210
rect 194 -211 195 -210
rect 195 -211 196 -210
rect 196 -211 197 -210
rect 197 -211 198 -210
rect 198 -211 199 -210
rect 199 -211 200 -210
rect 200 -211 201 -210
rect 201 -211 202 -210
rect 202 -211 203 -210
rect 203 -211 204 -210
rect 204 -211 205 -210
rect 205 -211 206 -210
rect 206 -211 207 -210
rect 207 -211 208 -210
rect 208 -211 209 -210
rect 209 -211 210 -210
rect 210 -211 211 -210
rect 211 -211 212 -210
rect 212 -211 213 -210
rect 213 -211 214 -210
rect 214 -211 215 -210
rect 215 -211 216 -210
rect 216 -211 217 -210
rect 217 -211 218 -210
rect 218 -211 219 -210
rect 219 -211 220 -210
rect 220 -211 221 -210
rect 221 -211 222 -210
rect 222 -211 223 -210
rect 223 -211 224 -210
rect 224 -211 225 -210
rect 225 -211 226 -210
rect 226 -211 227 -210
rect 227 -211 228 -210
rect 228 -211 229 -210
rect 229 -211 230 -210
rect 230 -211 231 -210
rect 231 -211 232 -210
rect 232 -211 233 -210
rect 233 -211 234 -210
rect 234 -211 235 -210
rect 235 -211 236 -210
rect 236 -211 237 -210
rect 237 -211 238 -210
rect 238 -211 239 -210
rect 239 -211 240 -210
rect 240 -211 241 -210
rect 241 -211 242 -210
rect 242 -211 243 -210
rect 243 -211 244 -210
rect 244 -211 245 -210
rect 245 -211 246 -210
rect 246 -211 247 -210
rect 247 -211 248 -210
rect 248 -211 249 -210
rect 249 -211 250 -210
rect 250 -211 251 -210
rect 251 -211 252 -210
rect 252 -211 253 -210
rect 253 -211 254 -210
rect 254 -211 255 -210
rect 255 -211 256 -210
rect 256 -211 257 -210
rect 257 -211 258 -210
rect 258 -211 259 -210
rect 259 -211 260 -210
rect 260 -211 261 -210
rect 261 -211 262 -210
rect 262 -211 263 -210
rect 263 -211 264 -210
rect 264 -211 265 -210
rect 265 -211 266 -210
rect 266 -211 267 -210
rect 267 -211 268 -210
rect 268 -211 269 -210
rect 269 -211 270 -210
rect 270 -211 271 -210
rect 271 -211 272 -210
rect 272 -211 273 -210
rect 273 -211 274 -210
rect 274 -211 275 -210
rect 275 -211 276 -210
rect 276 -211 277 -210
rect 277 -211 278 -210
rect 278 -211 279 -210
rect 279 -211 280 -210
rect 280 -211 281 -210
rect 281 -211 282 -210
rect 282 -211 283 -210
rect 283 -211 284 -210
rect 284 -211 285 -210
rect 285 -211 286 -210
rect 286 -211 287 -210
rect 287 -211 288 -210
rect 288 -211 289 -210
rect 289 -211 290 -210
rect 290 -211 291 -210
rect 291 -211 292 -210
rect 292 -211 293 -210
rect 293 -211 294 -210
rect 294 -211 295 -210
rect 295 -211 296 -210
rect 296 -211 297 -210
rect 297 -211 298 -210
rect 298 -211 299 -210
rect 299 -211 300 -210
rect 300 -211 301 -210
rect 301 -211 302 -210
rect 302 -211 303 -210
rect 303 -211 304 -210
rect 304 -211 305 -210
rect 305 -211 306 -210
rect 306 -211 307 -210
rect 307 -211 308 -210
rect 308 -211 309 -210
rect 309 -211 310 -210
rect 310 -211 311 -210
rect 311 -211 312 -210
rect 312 -211 313 -210
rect 313 -211 314 -210
rect 314 -211 315 -210
rect 315 -211 316 -210
rect 316 -211 317 -210
rect 317 -211 318 -210
rect 318 -211 319 -210
rect 319 -211 320 -210
rect 320 -211 321 -210
rect 321 -211 322 -210
rect 322 -211 323 -210
rect 323 -211 324 -210
rect 324 -211 325 -210
rect 325 -211 326 -210
rect 326 -211 327 -210
rect 327 -211 328 -210
rect 328 -211 329 -210
rect 329 -211 330 -210
rect 330 -211 331 -210
rect 331 -211 332 -210
rect 332 -211 333 -210
rect 333 -211 334 -210
rect 334 -211 335 -210
rect 335 -211 336 -210
rect 336 -211 337 -210
rect 337 -211 338 -210
rect 338 -211 339 -210
rect 339 -211 340 -210
rect 340 -211 341 -210
rect 341 -211 342 -210
rect 342 -211 343 -210
rect 343 -211 344 -210
rect 344 -211 345 -210
rect 345 -211 346 -210
rect 346 -211 347 -210
rect 347 -211 348 -210
rect 348 -211 349 -210
rect 349 -211 350 -210
rect 350 -211 351 -210
rect 351 -211 352 -210
rect 352 -211 353 -210
rect 353 -211 354 -210
rect 354 -211 355 -210
rect 355 -211 356 -210
rect 356 -211 357 -210
rect 357 -211 358 -210
rect 358 -211 359 -210
rect 359 -211 360 -210
rect 360 -211 361 -210
rect 361 -211 362 -210
rect 362 -211 363 -210
rect 363 -211 364 -210
rect 364 -211 365 -210
rect 365 -211 366 -210
rect 366 -211 367 -210
rect 367 -211 368 -210
rect 368 -211 369 -210
rect 369 -211 370 -210
rect 370 -211 371 -210
rect 371 -211 372 -210
rect 372 -211 373 -210
rect 373 -211 374 -210
rect 374 -211 375 -210
rect 375 -211 376 -210
rect 376 -211 377 -210
rect 377 -211 378 -210
rect 378 -211 379 -210
rect 379 -211 380 -210
rect 380 -211 381 -210
rect 381 -211 382 -210
rect 382 -211 383 -210
rect 383 -211 384 -210
rect 384 -211 385 -210
rect 385 -211 386 -210
rect 386 -211 387 -210
rect 387 -211 388 -210
rect 388 -211 389 -210
rect 389 -211 390 -210
rect 390 -211 391 -210
rect 391 -211 392 -210
rect 392 -211 393 -210
rect 393 -211 394 -210
rect 394 -211 395 -210
rect 395 -211 396 -210
rect 396 -211 397 -210
rect 397 -211 398 -210
rect 398 -211 399 -210
rect 399 -211 400 -210
rect 400 -211 401 -210
rect 401 -211 402 -210
rect 402 -211 403 -210
rect 403 -211 404 -210
rect 404 -211 405 -210
rect 405 -211 406 -210
rect 406 -211 407 -210
rect 407 -211 408 -210
rect 408 -211 409 -210
rect 409 -211 410 -210
rect 410 -211 411 -210
rect 411 -211 412 -210
rect 412 -211 413 -210
rect 413 -211 414 -210
rect 414 -211 415 -210
rect 415 -211 416 -210
rect 416 -211 417 -210
rect 417 -211 418 -210
rect 418 -211 419 -210
rect 419 -211 420 -210
rect 420 -211 421 -210
rect 421 -211 422 -210
rect 422 -211 423 -210
rect 423 -211 424 -210
rect 424 -211 425 -210
rect 425 -211 426 -210
rect 426 -211 427 -210
rect 427 -211 428 -210
rect 428 -211 429 -210
rect 429 -211 430 -210
rect 430 -211 431 -210
rect 431 -211 432 -210
rect 432 -211 433 -210
rect 433 -211 434 -210
rect 434 -211 435 -210
rect 435 -211 436 -210
rect 436 -211 437 -210
rect 437 -211 438 -210
rect 438 -211 439 -210
rect 439 -211 440 -210
rect 440 -211 441 -210
rect 441 -211 442 -210
rect 442 -211 443 -210
rect 443 -211 444 -210
rect 444 -211 445 -210
rect 445 -211 446 -210
rect 446 -211 447 -210
rect 447 -211 448 -210
rect 448 -211 449 -210
rect 449 -211 450 -210
rect 450 -211 451 -210
rect 451 -211 452 -210
rect 452 -211 453 -210
rect 453 -211 454 -210
rect 454 -211 455 -210
rect 455 -211 456 -210
rect 456 -211 457 -210
rect 457 -211 458 -210
rect 458 -211 459 -210
rect 459 -211 460 -210
rect 460 -211 461 -210
rect 461 -211 462 -210
rect 462 -211 463 -210
rect 463 -211 464 -210
rect 464 -211 465 -210
rect 465 -211 466 -210
rect 466 -211 467 -210
rect 467 -211 468 -210
rect 468 -211 469 -210
rect 469 -211 470 -210
rect 470 -211 471 -210
rect 471 -211 472 -210
rect 472 -211 473 -210
rect 473 -211 474 -210
rect 474 -211 475 -210
rect 475 -211 476 -210
rect 476 -211 477 -210
rect 477 -211 478 -210
rect 478 -211 479 -210
rect 479 -211 480 -210
rect 2 -212 3 -211
rect 3 -212 4 -211
rect 4 -212 5 -211
rect 5 -212 6 -211
rect 6 -212 7 -211
rect 7 -212 8 -211
rect 8 -212 9 -211
rect 9 -212 10 -211
rect 10 -212 11 -211
rect 11 -212 12 -211
rect 12 -212 13 -211
rect 13 -212 14 -211
rect 14 -212 15 -211
rect 15 -212 16 -211
rect 16 -212 17 -211
rect 17 -212 18 -211
rect 18 -212 19 -211
rect 19 -212 20 -211
rect 20 -212 21 -211
rect 21 -212 22 -211
rect 22 -212 23 -211
rect 23 -212 24 -211
rect 24 -212 25 -211
rect 25 -212 26 -211
rect 26 -212 27 -211
rect 27 -212 28 -211
rect 28 -212 29 -211
rect 29 -212 30 -211
rect 30 -212 31 -211
rect 31 -212 32 -211
rect 32 -212 33 -211
rect 33 -212 34 -211
rect 34 -212 35 -211
rect 35 -212 36 -211
rect 36 -212 37 -211
rect 37 -212 38 -211
rect 38 -212 39 -211
rect 39 -212 40 -211
rect 40 -212 41 -211
rect 41 -212 42 -211
rect 42 -212 43 -211
rect 43 -212 44 -211
rect 44 -212 45 -211
rect 45 -212 46 -211
rect 46 -212 47 -211
rect 47 -212 48 -211
rect 48 -212 49 -211
rect 49 -212 50 -211
rect 50 -212 51 -211
rect 51 -212 52 -211
rect 52 -212 53 -211
rect 53 -212 54 -211
rect 54 -212 55 -211
rect 55 -212 56 -211
rect 56 -212 57 -211
rect 57 -212 58 -211
rect 58 -212 59 -211
rect 59 -212 60 -211
rect 60 -212 61 -211
rect 61 -212 62 -211
rect 62 -212 63 -211
rect 63 -212 64 -211
rect 64 -212 65 -211
rect 65 -212 66 -211
rect 66 -212 67 -211
rect 67 -212 68 -211
rect 68 -212 69 -211
rect 69 -212 70 -211
rect 70 -212 71 -211
rect 71 -212 72 -211
rect 72 -212 73 -211
rect 73 -212 74 -211
rect 74 -212 75 -211
rect 75 -212 76 -211
rect 76 -212 77 -211
rect 77 -212 78 -211
rect 78 -212 79 -211
rect 79 -212 80 -211
rect 80 -212 81 -211
rect 81 -212 82 -211
rect 82 -212 83 -211
rect 83 -212 84 -211
rect 84 -212 85 -211
rect 85 -212 86 -211
rect 86 -212 87 -211
rect 87 -212 88 -211
rect 88 -212 89 -211
rect 89 -212 90 -211
rect 90 -212 91 -211
rect 91 -212 92 -211
rect 92 -212 93 -211
rect 93 -212 94 -211
rect 94 -212 95 -211
rect 95 -212 96 -211
rect 96 -212 97 -211
rect 97 -212 98 -211
rect 98 -212 99 -211
rect 99 -212 100 -211
rect 100 -212 101 -211
rect 101 -212 102 -211
rect 102 -212 103 -211
rect 103 -212 104 -211
rect 104 -212 105 -211
rect 105 -212 106 -211
rect 106 -212 107 -211
rect 107 -212 108 -211
rect 108 -212 109 -211
rect 109 -212 110 -211
rect 110 -212 111 -211
rect 111 -212 112 -211
rect 112 -212 113 -211
rect 113 -212 114 -211
rect 114 -212 115 -211
rect 115 -212 116 -211
rect 116 -212 117 -211
rect 117 -212 118 -211
rect 118 -212 119 -211
rect 119 -212 120 -211
rect 120 -212 121 -211
rect 121 -212 122 -211
rect 122 -212 123 -211
rect 123 -212 124 -211
rect 124 -212 125 -211
rect 125 -212 126 -211
rect 126 -212 127 -211
rect 127 -212 128 -211
rect 128 -212 129 -211
rect 129 -212 130 -211
rect 130 -212 131 -211
rect 131 -212 132 -211
rect 132 -212 133 -211
rect 133 -212 134 -211
rect 134 -212 135 -211
rect 135 -212 136 -211
rect 136 -212 137 -211
rect 137 -212 138 -211
rect 138 -212 139 -211
rect 139 -212 140 -211
rect 140 -212 141 -211
rect 141 -212 142 -211
rect 142 -212 143 -211
rect 143 -212 144 -211
rect 144 -212 145 -211
rect 145 -212 146 -211
rect 146 -212 147 -211
rect 147 -212 148 -211
rect 148 -212 149 -211
rect 149 -212 150 -211
rect 150 -212 151 -211
rect 151 -212 152 -211
rect 152 -212 153 -211
rect 153 -212 154 -211
rect 154 -212 155 -211
rect 155 -212 156 -211
rect 156 -212 157 -211
rect 157 -212 158 -211
rect 158 -212 159 -211
rect 159 -212 160 -211
rect 160 -212 161 -211
rect 161 -212 162 -211
rect 162 -212 163 -211
rect 163 -212 164 -211
rect 164 -212 165 -211
rect 165 -212 166 -211
rect 166 -212 167 -211
rect 167 -212 168 -211
rect 168 -212 169 -211
rect 169 -212 170 -211
rect 170 -212 171 -211
rect 171 -212 172 -211
rect 172 -212 173 -211
rect 173 -212 174 -211
rect 174 -212 175 -211
rect 175 -212 176 -211
rect 176 -212 177 -211
rect 177 -212 178 -211
rect 178 -212 179 -211
rect 179 -212 180 -211
rect 180 -212 181 -211
rect 181 -212 182 -211
rect 182 -212 183 -211
rect 183 -212 184 -211
rect 184 -212 185 -211
rect 185 -212 186 -211
rect 186 -212 187 -211
rect 187 -212 188 -211
rect 188 -212 189 -211
rect 189 -212 190 -211
rect 190 -212 191 -211
rect 191 -212 192 -211
rect 192 -212 193 -211
rect 193 -212 194 -211
rect 194 -212 195 -211
rect 195 -212 196 -211
rect 196 -212 197 -211
rect 197 -212 198 -211
rect 198 -212 199 -211
rect 199 -212 200 -211
rect 200 -212 201 -211
rect 201 -212 202 -211
rect 202 -212 203 -211
rect 203 -212 204 -211
rect 204 -212 205 -211
rect 205 -212 206 -211
rect 206 -212 207 -211
rect 207 -212 208 -211
rect 208 -212 209 -211
rect 209 -212 210 -211
rect 210 -212 211 -211
rect 211 -212 212 -211
rect 212 -212 213 -211
rect 213 -212 214 -211
rect 214 -212 215 -211
rect 215 -212 216 -211
rect 216 -212 217 -211
rect 217 -212 218 -211
rect 218 -212 219 -211
rect 219 -212 220 -211
rect 220 -212 221 -211
rect 221 -212 222 -211
rect 222 -212 223 -211
rect 223 -212 224 -211
rect 224 -212 225 -211
rect 225 -212 226 -211
rect 226 -212 227 -211
rect 227 -212 228 -211
rect 228 -212 229 -211
rect 229 -212 230 -211
rect 230 -212 231 -211
rect 231 -212 232 -211
rect 232 -212 233 -211
rect 233 -212 234 -211
rect 234 -212 235 -211
rect 235 -212 236 -211
rect 236 -212 237 -211
rect 237 -212 238 -211
rect 238 -212 239 -211
rect 239 -212 240 -211
rect 240 -212 241 -211
rect 241 -212 242 -211
rect 242 -212 243 -211
rect 243 -212 244 -211
rect 244 -212 245 -211
rect 245 -212 246 -211
rect 246 -212 247 -211
rect 247 -212 248 -211
rect 248 -212 249 -211
rect 249 -212 250 -211
rect 250 -212 251 -211
rect 251 -212 252 -211
rect 252 -212 253 -211
rect 253 -212 254 -211
rect 254 -212 255 -211
rect 255 -212 256 -211
rect 256 -212 257 -211
rect 257 -212 258 -211
rect 258 -212 259 -211
rect 259 -212 260 -211
rect 260 -212 261 -211
rect 261 -212 262 -211
rect 262 -212 263 -211
rect 263 -212 264 -211
rect 264 -212 265 -211
rect 265 -212 266 -211
rect 266 -212 267 -211
rect 267 -212 268 -211
rect 268 -212 269 -211
rect 269 -212 270 -211
rect 270 -212 271 -211
rect 271 -212 272 -211
rect 272 -212 273 -211
rect 273 -212 274 -211
rect 274 -212 275 -211
rect 275 -212 276 -211
rect 276 -212 277 -211
rect 277 -212 278 -211
rect 278 -212 279 -211
rect 279 -212 280 -211
rect 280 -212 281 -211
rect 281 -212 282 -211
rect 282 -212 283 -211
rect 283 -212 284 -211
rect 284 -212 285 -211
rect 285 -212 286 -211
rect 286 -212 287 -211
rect 287 -212 288 -211
rect 288 -212 289 -211
rect 289 -212 290 -211
rect 290 -212 291 -211
rect 291 -212 292 -211
rect 292 -212 293 -211
rect 293 -212 294 -211
rect 294 -212 295 -211
rect 295 -212 296 -211
rect 296 -212 297 -211
rect 297 -212 298 -211
rect 298 -212 299 -211
rect 299 -212 300 -211
rect 300 -212 301 -211
rect 301 -212 302 -211
rect 302 -212 303 -211
rect 303 -212 304 -211
rect 304 -212 305 -211
rect 305 -212 306 -211
rect 306 -212 307 -211
rect 307 -212 308 -211
rect 308 -212 309 -211
rect 309 -212 310 -211
rect 310 -212 311 -211
rect 311 -212 312 -211
rect 312 -212 313 -211
rect 313 -212 314 -211
rect 314 -212 315 -211
rect 315 -212 316 -211
rect 316 -212 317 -211
rect 317 -212 318 -211
rect 318 -212 319 -211
rect 319 -212 320 -211
rect 320 -212 321 -211
rect 321 -212 322 -211
rect 322 -212 323 -211
rect 323 -212 324 -211
rect 324 -212 325 -211
rect 325 -212 326 -211
rect 326 -212 327 -211
rect 327 -212 328 -211
rect 328 -212 329 -211
rect 329 -212 330 -211
rect 330 -212 331 -211
rect 331 -212 332 -211
rect 332 -212 333 -211
rect 333 -212 334 -211
rect 334 -212 335 -211
rect 335 -212 336 -211
rect 336 -212 337 -211
rect 337 -212 338 -211
rect 338 -212 339 -211
rect 339 -212 340 -211
rect 340 -212 341 -211
rect 341 -212 342 -211
rect 342 -212 343 -211
rect 343 -212 344 -211
rect 344 -212 345 -211
rect 345 -212 346 -211
rect 346 -212 347 -211
rect 347 -212 348 -211
rect 348 -212 349 -211
rect 349 -212 350 -211
rect 350 -212 351 -211
rect 351 -212 352 -211
rect 352 -212 353 -211
rect 353 -212 354 -211
rect 354 -212 355 -211
rect 355 -212 356 -211
rect 356 -212 357 -211
rect 357 -212 358 -211
rect 358 -212 359 -211
rect 359 -212 360 -211
rect 360 -212 361 -211
rect 361 -212 362 -211
rect 362 -212 363 -211
rect 363 -212 364 -211
rect 364 -212 365 -211
rect 365 -212 366 -211
rect 366 -212 367 -211
rect 367 -212 368 -211
rect 368 -212 369 -211
rect 369 -212 370 -211
rect 370 -212 371 -211
rect 371 -212 372 -211
rect 372 -212 373 -211
rect 373 -212 374 -211
rect 374 -212 375 -211
rect 375 -212 376 -211
rect 376 -212 377 -211
rect 377 -212 378 -211
rect 378 -212 379 -211
rect 379 -212 380 -211
rect 380 -212 381 -211
rect 381 -212 382 -211
rect 382 -212 383 -211
rect 383 -212 384 -211
rect 384 -212 385 -211
rect 385 -212 386 -211
rect 386 -212 387 -211
rect 387 -212 388 -211
rect 388 -212 389 -211
rect 389 -212 390 -211
rect 390 -212 391 -211
rect 391 -212 392 -211
rect 392 -212 393 -211
rect 393 -212 394 -211
rect 394 -212 395 -211
rect 395 -212 396 -211
rect 396 -212 397 -211
rect 397 -212 398 -211
rect 398 -212 399 -211
rect 399 -212 400 -211
rect 400 -212 401 -211
rect 401 -212 402 -211
rect 402 -212 403 -211
rect 403 -212 404 -211
rect 404 -212 405 -211
rect 405 -212 406 -211
rect 406 -212 407 -211
rect 407 -212 408 -211
rect 408 -212 409 -211
rect 409 -212 410 -211
rect 410 -212 411 -211
rect 411 -212 412 -211
rect 412 -212 413 -211
rect 413 -212 414 -211
rect 414 -212 415 -211
rect 415 -212 416 -211
rect 416 -212 417 -211
rect 417 -212 418 -211
rect 418 -212 419 -211
rect 419 -212 420 -211
rect 420 -212 421 -211
rect 421 -212 422 -211
rect 422 -212 423 -211
rect 423 -212 424 -211
rect 424 -212 425 -211
rect 425 -212 426 -211
rect 426 -212 427 -211
rect 427 -212 428 -211
rect 428 -212 429 -211
rect 429 -212 430 -211
rect 430 -212 431 -211
rect 431 -212 432 -211
rect 432 -212 433 -211
rect 433 -212 434 -211
rect 434 -212 435 -211
rect 435 -212 436 -211
rect 436 -212 437 -211
rect 437 -212 438 -211
rect 438 -212 439 -211
rect 439 -212 440 -211
rect 440 -212 441 -211
rect 441 -212 442 -211
rect 442 -212 443 -211
rect 443 -212 444 -211
rect 444 -212 445 -211
rect 445 -212 446 -211
rect 446 -212 447 -211
rect 447 -212 448 -211
rect 448 -212 449 -211
rect 449 -212 450 -211
rect 450 -212 451 -211
rect 451 -212 452 -211
rect 452 -212 453 -211
rect 453 -212 454 -211
rect 454 -212 455 -211
rect 455 -212 456 -211
rect 456 -212 457 -211
rect 457 -212 458 -211
rect 458 -212 459 -211
rect 459 -212 460 -211
rect 460 -212 461 -211
rect 461 -212 462 -211
rect 462 -212 463 -211
rect 463 -212 464 -211
rect 464 -212 465 -211
rect 465 -212 466 -211
rect 466 -212 467 -211
rect 467 -212 468 -211
rect 468 -212 469 -211
rect 469 -212 470 -211
rect 470 -212 471 -211
rect 471 -212 472 -211
rect 472 -212 473 -211
rect 473 -212 474 -211
rect 474 -212 475 -211
rect 475 -212 476 -211
rect 476 -212 477 -211
rect 477 -212 478 -211
rect 478 -212 479 -211
rect 479 -212 480 -211
rect 2 -235 3 -234
rect 3 -235 4 -234
rect 4 -235 5 -234
rect 5 -235 6 -234
rect 6 -235 7 -234
rect 7 -235 8 -234
rect 8 -235 9 -234
rect 9 -235 10 -234
rect 10 -235 11 -234
rect 11 -235 12 -234
rect 12 -235 13 -234
rect 13 -235 14 -234
rect 14 -235 15 -234
rect 15 -235 16 -234
rect 16 -235 17 -234
rect 17 -235 18 -234
rect 18 -235 19 -234
rect 19 -235 20 -234
rect 20 -235 21 -234
rect 21 -235 22 -234
rect 22 -235 23 -234
rect 23 -235 24 -234
rect 24 -235 25 -234
rect 25 -235 26 -234
rect 26 -235 27 -234
rect 27 -235 28 -234
rect 28 -235 29 -234
rect 29 -235 30 -234
rect 30 -235 31 -234
rect 31 -235 32 -234
rect 32 -235 33 -234
rect 33 -235 34 -234
rect 34 -235 35 -234
rect 35 -235 36 -234
rect 36 -235 37 -234
rect 37 -235 38 -234
rect 38 -235 39 -234
rect 39 -235 40 -234
rect 40 -235 41 -234
rect 41 -235 42 -234
rect 42 -235 43 -234
rect 43 -235 44 -234
rect 44 -235 45 -234
rect 45 -235 46 -234
rect 46 -235 47 -234
rect 47 -235 48 -234
rect 48 -235 49 -234
rect 49 -235 50 -234
rect 50 -235 51 -234
rect 51 -235 52 -234
rect 52 -235 53 -234
rect 53 -235 54 -234
rect 54 -235 55 -234
rect 55 -235 56 -234
rect 56 -235 57 -234
rect 57 -235 58 -234
rect 58 -235 59 -234
rect 59 -235 60 -234
rect 60 -235 61 -234
rect 61 -235 62 -234
rect 62 -235 63 -234
rect 63 -235 64 -234
rect 64 -235 65 -234
rect 65 -235 66 -234
rect 66 -235 67 -234
rect 67 -235 68 -234
rect 68 -235 69 -234
rect 69 -235 70 -234
rect 70 -235 71 -234
rect 71 -235 72 -234
rect 72 -235 73 -234
rect 73 -235 74 -234
rect 74 -235 75 -234
rect 75 -235 76 -234
rect 76 -235 77 -234
rect 77 -235 78 -234
rect 78 -235 79 -234
rect 79 -235 80 -234
rect 80 -235 81 -234
rect 81 -235 82 -234
rect 82 -235 83 -234
rect 83 -235 84 -234
rect 84 -235 85 -234
rect 85 -235 86 -234
rect 86 -235 87 -234
rect 87 -235 88 -234
rect 88 -235 89 -234
rect 89 -235 90 -234
rect 90 -235 91 -234
rect 91 -235 92 -234
rect 92 -235 93 -234
rect 93 -235 94 -234
rect 94 -235 95 -234
rect 95 -235 96 -234
rect 96 -235 97 -234
rect 97 -235 98 -234
rect 98 -235 99 -234
rect 99 -235 100 -234
rect 100 -235 101 -234
rect 101 -235 102 -234
rect 102 -235 103 -234
rect 103 -235 104 -234
rect 104 -235 105 -234
rect 105 -235 106 -234
rect 106 -235 107 -234
rect 107 -235 108 -234
rect 108 -235 109 -234
rect 109 -235 110 -234
rect 110 -235 111 -234
rect 111 -235 112 -234
rect 112 -235 113 -234
rect 113 -235 114 -234
rect 114 -235 115 -234
rect 115 -235 116 -234
rect 116 -235 117 -234
rect 117 -235 118 -234
rect 118 -235 119 -234
rect 119 -235 120 -234
rect 120 -235 121 -234
rect 121 -235 122 -234
rect 122 -235 123 -234
rect 123 -235 124 -234
rect 124 -235 125 -234
rect 125 -235 126 -234
rect 126 -235 127 -234
rect 127 -235 128 -234
rect 128 -235 129 -234
rect 129 -235 130 -234
rect 130 -235 131 -234
rect 131 -235 132 -234
rect 132 -235 133 -234
rect 133 -235 134 -234
rect 134 -235 135 -234
rect 135 -235 136 -234
rect 136 -235 137 -234
rect 137 -235 138 -234
rect 138 -235 139 -234
rect 139 -235 140 -234
rect 140 -235 141 -234
rect 141 -235 142 -234
rect 142 -235 143 -234
rect 143 -235 144 -234
rect 144 -235 145 -234
rect 145 -235 146 -234
rect 146 -235 147 -234
rect 147 -235 148 -234
rect 148 -235 149 -234
rect 149 -235 150 -234
rect 150 -235 151 -234
rect 151 -235 152 -234
rect 152 -235 153 -234
rect 153 -235 154 -234
rect 154 -235 155 -234
rect 155 -235 156 -234
rect 156 -235 157 -234
rect 157 -235 158 -234
rect 158 -235 159 -234
rect 159 -235 160 -234
rect 160 -235 161 -234
rect 161 -235 162 -234
rect 162 -235 163 -234
rect 163 -235 164 -234
rect 164 -235 165 -234
rect 165 -235 166 -234
rect 166 -235 167 -234
rect 167 -235 168 -234
rect 168 -235 169 -234
rect 169 -235 170 -234
rect 170 -235 171 -234
rect 171 -235 172 -234
rect 172 -235 173 -234
rect 173 -235 174 -234
rect 174 -235 175 -234
rect 175 -235 176 -234
rect 176 -235 177 -234
rect 177 -235 178 -234
rect 178 -235 179 -234
rect 179 -235 180 -234
rect 180 -235 181 -234
rect 181 -235 182 -234
rect 182 -235 183 -234
rect 183 -235 184 -234
rect 184 -235 185 -234
rect 185 -235 186 -234
rect 186 -235 187 -234
rect 187 -235 188 -234
rect 188 -235 189 -234
rect 189 -235 190 -234
rect 190 -235 191 -234
rect 191 -235 192 -234
rect 192 -235 193 -234
rect 193 -235 194 -234
rect 194 -235 195 -234
rect 195 -235 196 -234
rect 196 -235 197 -234
rect 197 -235 198 -234
rect 198 -235 199 -234
rect 199 -235 200 -234
rect 200 -235 201 -234
rect 201 -235 202 -234
rect 202 -235 203 -234
rect 203 -235 204 -234
rect 204 -235 205 -234
rect 205 -235 206 -234
rect 206 -235 207 -234
rect 207 -235 208 -234
rect 208 -235 209 -234
rect 209 -235 210 -234
rect 210 -235 211 -234
rect 211 -235 212 -234
rect 212 -235 213 -234
rect 213 -235 214 -234
rect 214 -235 215 -234
rect 215 -235 216 -234
rect 216 -235 217 -234
rect 217 -235 218 -234
rect 218 -235 219 -234
rect 219 -235 220 -234
rect 220 -235 221 -234
rect 221 -235 222 -234
rect 222 -235 223 -234
rect 223 -235 224 -234
rect 224 -235 225 -234
rect 225 -235 226 -234
rect 226 -235 227 -234
rect 227 -235 228 -234
rect 228 -235 229 -234
rect 229 -235 230 -234
rect 230 -235 231 -234
rect 231 -235 232 -234
rect 232 -235 233 -234
rect 233 -235 234 -234
rect 234 -235 235 -234
rect 235 -235 236 -234
rect 236 -235 237 -234
rect 237 -235 238 -234
rect 238 -235 239 -234
rect 239 -235 240 -234
rect 240 -235 241 -234
rect 241 -235 242 -234
rect 242 -235 243 -234
rect 243 -235 244 -234
rect 244 -235 245 -234
rect 245 -235 246 -234
rect 246 -235 247 -234
rect 247 -235 248 -234
rect 248 -235 249 -234
rect 249 -235 250 -234
rect 250 -235 251 -234
rect 251 -235 252 -234
rect 252 -235 253 -234
rect 253 -235 254 -234
rect 254 -235 255 -234
rect 255 -235 256 -234
rect 256 -235 257 -234
rect 257 -235 258 -234
rect 258 -235 259 -234
rect 259 -235 260 -234
rect 260 -235 261 -234
rect 261 -235 262 -234
rect 262 -235 263 -234
rect 263 -235 264 -234
rect 264 -235 265 -234
rect 265 -235 266 -234
rect 266 -235 267 -234
rect 267 -235 268 -234
rect 268 -235 269 -234
rect 269 -235 270 -234
rect 270 -235 271 -234
rect 271 -235 272 -234
rect 272 -235 273 -234
rect 273 -235 274 -234
rect 274 -235 275 -234
rect 275 -235 276 -234
rect 276 -235 277 -234
rect 277 -235 278 -234
rect 278 -235 279 -234
rect 279 -235 280 -234
rect 280 -235 281 -234
rect 281 -235 282 -234
rect 282 -235 283 -234
rect 283 -235 284 -234
rect 284 -235 285 -234
rect 285 -235 286 -234
rect 286 -235 287 -234
rect 287 -235 288 -234
rect 288 -235 289 -234
rect 289 -235 290 -234
rect 290 -235 291 -234
rect 291 -235 292 -234
rect 292 -235 293 -234
rect 293 -235 294 -234
rect 294 -235 295 -234
rect 295 -235 296 -234
rect 296 -235 297 -234
rect 297 -235 298 -234
rect 298 -235 299 -234
rect 299 -235 300 -234
rect 300 -235 301 -234
rect 301 -235 302 -234
rect 302 -235 303 -234
rect 303 -235 304 -234
rect 304 -235 305 -234
rect 305 -235 306 -234
rect 306 -235 307 -234
rect 307 -235 308 -234
rect 308 -235 309 -234
rect 309 -235 310 -234
rect 310 -235 311 -234
rect 311 -235 312 -234
rect 312 -235 313 -234
rect 313 -235 314 -234
rect 314 -235 315 -234
rect 315 -235 316 -234
rect 316 -235 317 -234
rect 317 -235 318 -234
rect 318 -235 319 -234
rect 319 -235 320 -234
rect 320 -235 321 -234
rect 321 -235 322 -234
rect 322 -235 323 -234
rect 323 -235 324 -234
rect 324 -235 325 -234
rect 325 -235 326 -234
rect 326 -235 327 -234
rect 327 -235 328 -234
rect 328 -235 329 -234
rect 329 -235 330 -234
rect 330 -235 331 -234
rect 331 -235 332 -234
rect 332 -235 333 -234
rect 333 -235 334 -234
rect 334 -235 335 -234
rect 335 -235 336 -234
rect 336 -235 337 -234
rect 337 -235 338 -234
rect 338 -235 339 -234
rect 339 -235 340 -234
rect 340 -235 341 -234
rect 341 -235 342 -234
rect 342 -235 343 -234
rect 343 -235 344 -234
rect 344 -235 345 -234
rect 345 -235 346 -234
rect 346 -235 347 -234
rect 347 -235 348 -234
rect 348 -235 349 -234
rect 349 -235 350 -234
rect 350 -235 351 -234
rect 351 -235 352 -234
rect 352 -235 353 -234
rect 353 -235 354 -234
rect 354 -235 355 -234
rect 355 -235 356 -234
rect 356 -235 357 -234
rect 357 -235 358 -234
rect 358 -235 359 -234
rect 359 -235 360 -234
rect 360 -235 361 -234
rect 361 -235 362 -234
rect 362 -235 363 -234
rect 363 -235 364 -234
rect 364 -235 365 -234
rect 365 -235 366 -234
rect 366 -235 367 -234
rect 367 -235 368 -234
rect 368 -235 369 -234
rect 369 -235 370 -234
rect 370 -235 371 -234
rect 371 -235 372 -234
rect 372 -235 373 -234
rect 373 -235 374 -234
rect 374 -235 375 -234
rect 375 -235 376 -234
rect 376 -235 377 -234
rect 377 -235 378 -234
rect 378 -235 379 -234
rect 379 -235 380 -234
rect 380 -235 381 -234
rect 381 -235 382 -234
rect 382 -235 383 -234
rect 383 -235 384 -234
rect 384 -235 385 -234
rect 385 -235 386 -234
rect 386 -235 387 -234
rect 387 -235 388 -234
rect 388 -235 389 -234
rect 389 -235 390 -234
rect 390 -235 391 -234
rect 391 -235 392 -234
rect 392 -235 393 -234
rect 393 -235 394 -234
rect 394 -235 395 -234
rect 395 -235 396 -234
rect 396 -235 397 -234
rect 397 -235 398 -234
rect 398 -235 399 -234
rect 399 -235 400 -234
rect 400 -235 401 -234
rect 401 -235 402 -234
rect 402 -235 403 -234
rect 403 -235 404 -234
rect 404 -235 405 -234
rect 405 -235 406 -234
rect 406 -235 407 -234
rect 407 -235 408 -234
rect 408 -235 409 -234
rect 409 -235 410 -234
rect 410 -235 411 -234
rect 411 -235 412 -234
rect 412 -235 413 -234
rect 413 -235 414 -234
rect 414 -235 415 -234
rect 415 -235 416 -234
rect 416 -235 417 -234
rect 417 -235 418 -234
rect 418 -235 419 -234
rect 419 -235 420 -234
rect 420 -235 421 -234
rect 421 -235 422 -234
rect 422 -235 423 -234
rect 423 -235 424 -234
rect 424 -235 425 -234
rect 425 -235 426 -234
rect 426 -235 427 -234
rect 427 -235 428 -234
rect 428 -235 429 -234
rect 429 -235 430 -234
rect 430 -235 431 -234
rect 431 -235 432 -234
rect 432 -235 433 -234
rect 433 -235 434 -234
rect 434 -235 435 -234
rect 435 -235 436 -234
rect 436 -235 437 -234
rect 437 -235 438 -234
rect 438 -235 439 -234
rect 439 -235 440 -234
rect 440 -235 441 -234
rect 441 -235 442 -234
rect 442 -235 443 -234
rect 443 -235 444 -234
rect 444 -235 445 -234
rect 445 -235 446 -234
rect 446 -235 447 -234
rect 447 -235 448 -234
rect 448 -235 449 -234
rect 449 -235 450 -234
rect 450 -235 451 -234
rect 451 -235 452 -234
rect 452 -235 453 -234
rect 453 -235 454 -234
rect 454 -235 455 -234
rect 455 -235 456 -234
rect 456 -235 457 -234
rect 457 -235 458 -234
rect 458 -235 459 -234
rect 459 -235 460 -234
rect 460 -235 461 -234
rect 461 -235 462 -234
rect 462 -235 463 -234
rect 463 -235 464 -234
rect 464 -235 465 -234
rect 465 -235 466 -234
rect 466 -235 467 -234
rect 467 -235 468 -234
rect 468 -235 469 -234
rect 469 -235 470 -234
rect 470 -235 471 -234
rect 471 -235 472 -234
rect 472 -235 473 -234
rect 473 -235 474 -234
rect 474 -235 475 -234
rect 475 -235 476 -234
rect 476 -235 477 -234
rect 477 -235 478 -234
rect 478 -235 479 -234
rect 479 -235 480 -234
rect 2 -236 3 -235
rect 3 -236 4 -235
rect 4 -236 5 -235
rect 5 -236 6 -235
rect 6 -236 7 -235
rect 7 -236 8 -235
rect 8 -236 9 -235
rect 9 -236 10 -235
rect 10 -236 11 -235
rect 11 -236 12 -235
rect 12 -236 13 -235
rect 13 -236 14 -235
rect 14 -236 15 -235
rect 15 -236 16 -235
rect 16 -236 17 -235
rect 17 -236 18 -235
rect 18 -236 19 -235
rect 19 -236 20 -235
rect 20 -236 21 -235
rect 21 -236 22 -235
rect 22 -236 23 -235
rect 23 -236 24 -235
rect 24 -236 25 -235
rect 25 -236 26 -235
rect 26 -236 27 -235
rect 27 -236 28 -235
rect 28 -236 29 -235
rect 29 -236 30 -235
rect 30 -236 31 -235
rect 31 -236 32 -235
rect 32 -236 33 -235
rect 33 -236 34 -235
rect 34 -236 35 -235
rect 35 -236 36 -235
rect 36 -236 37 -235
rect 37 -236 38 -235
rect 38 -236 39 -235
rect 39 -236 40 -235
rect 40 -236 41 -235
rect 41 -236 42 -235
rect 42 -236 43 -235
rect 43 -236 44 -235
rect 44 -236 45 -235
rect 45 -236 46 -235
rect 46 -236 47 -235
rect 47 -236 48 -235
rect 48 -236 49 -235
rect 49 -236 50 -235
rect 50 -236 51 -235
rect 51 -236 52 -235
rect 52 -236 53 -235
rect 53 -236 54 -235
rect 54 -236 55 -235
rect 55 -236 56 -235
rect 56 -236 57 -235
rect 57 -236 58 -235
rect 58 -236 59 -235
rect 59 -236 60 -235
rect 60 -236 61 -235
rect 61 -236 62 -235
rect 62 -236 63 -235
rect 63 -236 64 -235
rect 64 -236 65 -235
rect 65 -236 66 -235
rect 66 -236 67 -235
rect 67 -236 68 -235
rect 68 -236 69 -235
rect 69 -236 70 -235
rect 70 -236 71 -235
rect 71 -236 72 -235
rect 72 -236 73 -235
rect 73 -236 74 -235
rect 74 -236 75 -235
rect 75 -236 76 -235
rect 76 -236 77 -235
rect 77 -236 78 -235
rect 78 -236 79 -235
rect 79 -236 80 -235
rect 80 -236 81 -235
rect 81 -236 82 -235
rect 82 -236 83 -235
rect 83 -236 84 -235
rect 84 -236 85 -235
rect 85 -236 86 -235
rect 86 -236 87 -235
rect 87 -236 88 -235
rect 88 -236 89 -235
rect 89 -236 90 -235
rect 90 -236 91 -235
rect 91 -236 92 -235
rect 92 -236 93 -235
rect 93 -236 94 -235
rect 94 -236 95 -235
rect 95 -236 96 -235
rect 96 -236 97 -235
rect 97 -236 98 -235
rect 98 -236 99 -235
rect 99 -236 100 -235
rect 100 -236 101 -235
rect 101 -236 102 -235
rect 102 -236 103 -235
rect 103 -236 104 -235
rect 104 -236 105 -235
rect 105 -236 106 -235
rect 106 -236 107 -235
rect 107 -236 108 -235
rect 108 -236 109 -235
rect 109 -236 110 -235
rect 110 -236 111 -235
rect 111 -236 112 -235
rect 112 -236 113 -235
rect 113 -236 114 -235
rect 114 -236 115 -235
rect 115 -236 116 -235
rect 116 -236 117 -235
rect 117 -236 118 -235
rect 118 -236 119 -235
rect 119 -236 120 -235
rect 120 -236 121 -235
rect 121 -236 122 -235
rect 122 -236 123 -235
rect 123 -236 124 -235
rect 124 -236 125 -235
rect 125 -236 126 -235
rect 126 -236 127 -235
rect 127 -236 128 -235
rect 128 -236 129 -235
rect 129 -236 130 -235
rect 130 -236 131 -235
rect 131 -236 132 -235
rect 132 -236 133 -235
rect 133 -236 134 -235
rect 134 -236 135 -235
rect 135 -236 136 -235
rect 136 -236 137 -235
rect 137 -236 138 -235
rect 138 -236 139 -235
rect 139 -236 140 -235
rect 140 -236 141 -235
rect 141 -236 142 -235
rect 142 -236 143 -235
rect 143 -236 144 -235
rect 144 -236 145 -235
rect 145 -236 146 -235
rect 146 -236 147 -235
rect 147 -236 148 -235
rect 148 -236 149 -235
rect 149 -236 150 -235
rect 150 -236 151 -235
rect 151 -236 152 -235
rect 152 -236 153 -235
rect 153 -236 154 -235
rect 154 -236 155 -235
rect 155 -236 156 -235
rect 156 -236 157 -235
rect 157 -236 158 -235
rect 158 -236 159 -235
rect 159 -236 160 -235
rect 160 -236 161 -235
rect 161 -236 162 -235
rect 162 -236 163 -235
rect 163 -236 164 -235
rect 164 -236 165 -235
rect 165 -236 166 -235
rect 166 -236 167 -235
rect 167 -236 168 -235
rect 168 -236 169 -235
rect 169 -236 170 -235
rect 170 -236 171 -235
rect 171 -236 172 -235
rect 172 -236 173 -235
rect 173 -236 174 -235
rect 174 -236 175 -235
rect 175 -236 176 -235
rect 176 -236 177 -235
rect 177 -236 178 -235
rect 178 -236 179 -235
rect 179 -236 180 -235
rect 180 -236 181 -235
rect 181 -236 182 -235
rect 182 -236 183 -235
rect 183 -236 184 -235
rect 184 -236 185 -235
rect 185 -236 186 -235
rect 186 -236 187 -235
rect 187 -236 188 -235
rect 188 -236 189 -235
rect 189 -236 190 -235
rect 190 -236 191 -235
rect 191 -236 192 -235
rect 192 -236 193 -235
rect 193 -236 194 -235
rect 194 -236 195 -235
rect 195 -236 196 -235
rect 196 -236 197 -235
rect 197 -236 198 -235
rect 198 -236 199 -235
rect 199 -236 200 -235
rect 200 -236 201 -235
rect 201 -236 202 -235
rect 202 -236 203 -235
rect 203 -236 204 -235
rect 204 -236 205 -235
rect 205 -236 206 -235
rect 206 -236 207 -235
rect 207 -236 208 -235
rect 208 -236 209 -235
rect 209 -236 210 -235
rect 210 -236 211 -235
rect 211 -236 212 -235
rect 212 -236 213 -235
rect 213 -236 214 -235
rect 214 -236 215 -235
rect 215 -236 216 -235
rect 216 -236 217 -235
rect 217 -236 218 -235
rect 218 -236 219 -235
rect 219 -236 220 -235
rect 220 -236 221 -235
rect 221 -236 222 -235
rect 222 -236 223 -235
rect 223 -236 224 -235
rect 224 -236 225 -235
rect 225 -236 226 -235
rect 226 -236 227 -235
rect 227 -236 228 -235
rect 228 -236 229 -235
rect 229 -236 230 -235
rect 230 -236 231 -235
rect 231 -236 232 -235
rect 232 -236 233 -235
rect 233 -236 234 -235
rect 234 -236 235 -235
rect 235 -236 236 -235
rect 236 -236 237 -235
rect 237 -236 238 -235
rect 238 -236 239 -235
rect 239 -236 240 -235
rect 240 -236 241 -235
rect 241 -236 242 -235
rect 242 -236 243 -235
rect 243 -236 244 -235
rect 244 -236 245 -235
rect 245 -236 246 -235
rect 246 -236 247 -235
rect 247 -236 248 -235
rect 248 -236 249 -235
rect 249 -236 250 -235
rect 250 -236 251 -235
rect 251 -236 252 -235
rect 252 -236 253 -235
rect 253 -236 254 -235
rect 254 -236 255 -235
rect 255 -236 256 -235
rect 256 -236 257 -235
rect 257 -236 258 -235
rect 258 -236 259 -235
rect 259 -236 260 -235
rect 260 -236 261 -235
rect 261 -236 262 -235
rect 262 -236 263 -235
rect 263 -236 264 -235
rect 264 -236 265 -235
rect 265 -236 266 -235
rect 266 -236 267 -235
rect 267 -236 268 -235
rect 268 -236 269 -235
rect 269 -236 270 -235
rect 270 -236 271 -235
rect 271 -236 272 -235
rect 272 -236 273 -235
rect 273 -236 274 -235
rect 274 -236 275 -235
rect 275 -236 276 -235
rect 276 -236 277 -235
rect 277 -236 278 -235
rect 278 -236 279 -235
rect 279 -236 280 -235
rect 280 -236 281 -235
rect 281 -236 282 -235
rect 282 -236 283 -235
rect 283 -236 284 -235
rect 284 -236 285 -235
rect 285 -236 286 -235
rect 286 -236 287 -235
rect 287 -236 288 -235
rect 288 -236 289 -235
rect 289 -236 290 -235
rect 290 -236 291 -235
rect 291 -236 292 -235
rect 292 -236 293 -235
rect 293 -236 294 -235
rect 294 -236 295 -235
rect 295 -236 296 -235
rect 296 -236 297 -235
rect 297 -236 298 -235
rect 298 -236 299 -235
rect 299 -236 300 -235
rect 300 -236 301 -235
rect 301 -236 302 -235
rect 302 -236 303 -235
rect 303 -236 304 -235
rect 304 -236 305 -235
rect 305 -236 306 -235
rect 306 -236 307 -235
rect 307 -236 308 -235
rect 308 -236 309 -235
rect 309 -236 310 -235
rect 310 -236 311 -235
rect 311 -236 312 -235
rect 312 -236 313 -235
rect 313 -236 314 -235
rect 314 -236 315 -235
rect 315 -236 316 -235
rect 316 -236 317 -235
rect 317 -236 318 -235
rect 318 -236 319 -235
rect 319 -236 320 -235
rect 320 -236 321 -235
rect 321 -236 322 -235
rect 322 -236 323 -235
rect 323 -236 324 -235
rect 324 -236 325 -235
rect 325 -236 326 -235
rect 326 -236 327 -235
rect 327 -236 328 -235
rect 328 -236 329 -235
rect 329 -236 330 -235
rect 330 -236 331 -235
rect 331 -236 332 -235
rect 332 -236 333 -235
rect 333 -236 334 -235
rect 334 -236 335 -235
rect 335 -236 336 -235
rect 336 -236 337 -235
rect 337 -236 338 -235
rect 338 -236 339 -235
rect 339 -236 340 -235
rect 340 -236 341 -235
rect 341 -236 342 -235
rect 342 -236 343 -235
rect 343 -236 344 -235
rect 344 -236 345 -235
rect 345 -236 346 -235
rect 346 -236 347 -235
rect 347 -236 348 -235
rect 348 -236 349 -235
rect 349 -236 350 -235
rect 350 -236 351 -235
rect 351 -236 352 -235
rect 352 -236 353 -235
rect 353 -236 354 -235
rect 354 -236 355 -235
rect 355 -236 356 -235
rect 356 -236 357 -235
rect 357 -236 358 -235
rect 358 -236 359 -235
rect 359 -236 360 -235
rect 360 -236 361 -235
rect 361 -236 362 -235
rect 362 -236 363 -235
rect 363 -236 364 -235
rect 364 -236 365 -235
rect 365 -236 366 -235
rect 366 -236 367 -235
rect 367 -236 368 -235
rect 368 -236 369 -235
rect 369 -236 370 -235
rect 370 -236 371 -235
rect 371 -236 372 -235
rect 372 -236 373 -235
rect 373 -236 374 -235
rect 374 -236 375 -235
rect 375 -236 376 -235
rect 376 -236 377 -235
rect 377 -236 378 -235
rect 378 -236 379 -235
rect 379 -236 380 -235
rect 380 -236 381 -235
rect 381 -236 382 -235
rect 382 -236 383 -235
rect 383 -236 384 -235
rect 384 -236 385 -235
rect 385 -236 386 -235
rect 386 -236 387 -235
rect 387 -236 388 -235
rect 388 -236 389 -235
rect 389 -236 390 -235
rect 390 -236 391 -235
rect 391 -236 392 -235
rect 392 -236 393 -235
rect 393 -236 394 -235
rect 394 -236 395 -235
rect 395 -236 396 -235
rect 396 -236 397 -235
rect 397 -236 398 -235
rect 398 -236 399 -235
rect 399 -236 400 -235
rect 400 -236 401 -235
rect 401 -236 402 -235
rect 402 -236 403 -235
rect 403 -236 404 -235
rect 404 -236 405 -235
rect 405 -236 406 -235
rect 406 -236 407 -235
rect 407 -236 408 -235
rect 408 -236 409 -235
rect 409 -236 410 -235
rect 410 -236 411 -235
rect 411 -236 412 -235
rect 412 -236 413 -235
rect 413 -236 414 -235
rect 414 -236 415 -235
rect 415 -236 416 -235
rect 416 -236 417 -235
rect 417 -236 418 -235
rect 418 -236 419 -235
rect 419 -236 420 -235
rect 420 -236 421 -235
rect 421 -236 422 -235
rect 422 -236 423 -235
rect 423 -236 424 -235
rect 424 -236 425 -235
rect 425 -236 426 -235
rect 426 -236 427 -235
rect 427 -236 428 -235
rect 428 -236 429 -235
rect 429 -236 430 -235
rect 430 -236 431 -235
rect 431 -236 432 -235
rect 432 -236 433 -235
rect 433 -236 434 -235
rect 434 -236 435 -235
rect 435 -236 436 -235
rect 436 -236 437 -235
rect 437 -236 438 -235
rect 438 -236 439 -235
rect 439 -236 440 -235
rect 440 -236 441 -235
rect 441 -236 442 -235
rect 442 -236 443 -235
rect 443 -236 444 -235
rect 444 -236 445 -235
rect 445 -236 446 -235
rect 446 -236 447 -235
rect 447 -236 448 -235
rect 448 -236 449 -235
rect 449 -236 450 -235
rect 450 -236 451 -235
rect 451 -236 452 -235
rect 452 -236 453 -235
rect 453 -236 454 -235
rect 454 -236 455 -235
rect 455 -236 456 -235
rect 456 -236 457 -235
rect 457 -236 458 -235
rect 458 -236 459 -235
rect 459 -236 460 -235
rect 460 -236 461 -235
rect 461 -236 462 -235
rect 462 -236 463 -235
rect 463 -236 464 -235
rect 464 -236 465 -235
rect 465 -236 466 -235
rect 466 -236 467 -235
rect 467 -236 468 -235
rect 468 -236 469 -235
rect 469 -236 470 -235
rect 470 -236 471 -235
rect 471 -236 472 -235
rect 472 -236 473 -235
rect 473 -236 474 -235
rect 474 -236 475 -235
rect 475 -236 476 -235
rect 476 -236 477 -235
rect 477 -236 478 -235
rect 478 -236 479 -235
rect 479 -236 480 -235
rect 2 -237 3 -236
rect 3 -237 4 -236
rect 4 -237 5 -236
rect 5 -237 6 -236
rect 6 -237 7 -236
rect 7 -237 8 -236
rect 8 -237 9 -236
rect 9 -237 10 -236
rect 10 -237 11 -236
rect 11 -237 12 -236
rect 12 -237 13 -236
rect 13 -237 14 -236
rect 14 -237 15 -236
rect 15 -237 16 -236
rect 16 -237 17 -236
rect 17 -237 18 -236
rect 18 -237 19 -236
rect 19 -237 20 -236
rect 20 -237 21 -236
rect 21 -237 22 -236
rect 22 -237 23 -236
rect 23 -237 24 -236
rect 24 -237 25 -236
rect 25 -237 26 -236
rect 26 -237 27 -236
rect 27 -237 28 -236
rect 28 -237 29 -236
rect 29 -237 30 -236
rect 30 -237 31 -236
rect 31 -237 32 -236
rect 32 -237 33 -236
rect 33 -237 34 -236
rect 34 -237 35 -236
rect 35 -237 36 -236
rect 36 -237 37 -236
rect 37 -237 38 -236
rect 38 -237 39 -236
rect 39 -237 40 -236
rect 40 -237 41 -236
rect 41 -237 42 -236
rect 42 -237 43 -236
rect 43 -237 44 -236
rect 44 -237 45 -236
rect 45 -237 46 -236
rect 46 -237 47 -236
rect 47 -237 48 -236
rect 48 -237 49 -236
rect 49 -237 50 -236
rect 50 -237 51 -236
rect 51 -237 52 -236
rect 52 -237 53 -236
rect 53 -237 54 -236
rect 54 -237 55 -236
rect 55 -237 56 -236
rect 56 -237 57 -236
rect 57 -237 58 -236
rect 58 -237 59 -236
rect 59 -237 60 -236
rect 60 -237 61 -236
rect 61 -237 62 -236
rect 62 -237 63 -236
rect 63 -237 64 -236
rect 64 -237 65 -236
rect 65 -237 66 -236
rect 66 -237 67 -236
rect 67 -237 68 -236
rect 68 -237 69 -236
rect 69 -237 70 -236
rect 70 -237 71 -236
rect 71 -237 72 -236
rect 72 -237 73 -236
rect 73 -237 74 -236
rect 74 -237 75 -236
rect 75 -237 76 -236
rect 76 -237 77 -236
rect 77 -237 78 -236
rect 78 -237 79 -236
rect 79 -237 80 -236
rect 80 -237 81 -236
rect 81 -237 82 -236
rect 82 -237 83 -236
rect 83 -237 84 -236
rect 84 -237 85 -236
rect 85 -237 86 -236
rect 86 -237 87 -236
rect 87 -237 88 -236
rect 88 -237 89 -236
rect 89 -237 90 -236
rect 90 -237 91 -236
rect 91 -237 92 -236
rect 92 -237 93 -236
rect 93 -237 94 -236
rect 94 -237 95 -236
rect 95 -237 96 -236
rect 96 -237 97 -236
rect 97 -237 98 -236
rect 98 -237 99 -236
rect 99 -237 100 -236
rect 100 -237 101 -236
rect 101 -237 102 -236
rect 102 -237 103 -236
rect 103 -237 104 -236
rect 104 -237 105 -236
rect 105 -237 106 -236
rect 106 -237 107 -236
rect 107 -237 108 -236
rect 108 -237 109 -236
rect 109 -237 110 -236
rect 110 -237 111 -236
rect 111 -237 112 -236
rect 112 -237 113 -236
rect 113 -237 114 -236
rect 114 -237 115 -236
rect 115 -237 116 -236
rect 116 -237 117 -236
rect 117 -237 118 -236
rect 118 -237 119 -236
rect 119 -237 120 -236
rect 120 -237 121 -236
rect 121 -237 122 -236
rect 122 -237 123 -236
rect 123 -237 124 -236
rect 124 -237 125 -236
rect 125 -237 126 -236
rect 126 -237 127 -236
rect 127 -237 128 -236
rect 128 -237 129 -236
rect 129 -237 130 -236
rect 130 -237 131 -236
rect 131 -237 132 -236
rect 132 -237 133 -236
rect 133 -237 134 -236
rect 134 -237 135 -236
rect 135 -237 136 -236
rect 136 -237 137 -236
rect 137 -237 138 -236
rect 138 -237 139 -236
rect 139 -237 140 -236
rect 140 -237 141 -236
rect 141 -237 142 -236
rect 142 -237 143 -236
rect 143 -237 144 -236
rect 144 -237 145 -236
rect 145 -237 146 -236
rect 146 -237 147 -236
rect 147 -237 148 -236
rect 148 -237 149 -236
rect 149 -237 150 -236
rect 150 -237 151 -236
rect 151 -237 152 -236
rect 152 -237 153 -236
rect 153 -237 154 -236
rect 154 -237 155 -236
rect 155 -237 156 -236
rect 156 -237 157 -236
rect 157 -237 158 -236
rect 158 -237 159 -236
rect 159 -237 160 -236
rect 160 -237 161 -236
rect 161 -237 162 -236
rect 162 -237 163 -236
rect 163 -237 164 -236
rect 164 -237 165 -236
rect 165 -237 166 -236
rect 166 -237 167 -236
rect 167 -237 168 -236
rect 168 -237 169 -236
rect 169 -237 170 -236
rect 170 -237 171 -236
rect 171 -237 172 -236
rect 172 -237 173 -236
rect 173 -237 174 -236
rect 174 -237 175 -236
rect 175 -237 176 -236
rect 176 -237 177 -236
rect 177 -237 178 -236
rect 178 -237 179 -236
rect 179 -237 180 -236
rect 180 -237 181 -236
rect 181 -237 182 -236
rect 182 -237 183 -236
rect 183 -237 184 -236
rect 184 -237 185 -236
rect 185 -237 186 -236
rect 186 -237 187 -236
rect 187 -237 188 -236
rect 188 -237 189 -236
rect 189 -237 190 -236
rect 190 -237 191 -236
rect 191 -237 192 -236
rect 192 -237 193 -236
rect 193 -237 194 -236
rect 194 -237 195 -236
rect 195 -237 196 -236
rect 196 -237 197 -236
rect 197 -237 198 -236
rect 198 -237 199 -236
rect 199 -237 200 -236
rect 200 -237 201 -236
rect 201 -237 202 -236
rect 202 -237 203 -236
rect 203 -237 204 -236
rect 204 -237 205 -236
rect 205 -237 206 -236
rect 206 -237 207 -236
rect 207 -237 208 -236
rect 208 -237 209 -236
rect 209 -237 210 -236
rect 210 -237 211 -236
rect 211 -237 212 -236
rect 212 -237 213 -236
rect 213 -237 214 -236
rect 214 -237 215 -236
rect 215 -237 216 -236
rect 216 -237 217 -236
rect 217 -237 218 -236
rect 218 -237 219 -236
rect 219 -237 220 -236
rect 220 -237 221 -236
rect 221 -237 222 -236
rect 222 -237 223 -236
rect 223 -237 224 -236
rect 224 -237 225 -236
rect 225 -237 226 -236
rect 226 -237 227 -236
rect 227 -237 228 -236
rect 228 -237 229 -236
rect 229 -237 230 -236
rect 230 -237 231 -236
rect 231 -237 232 -236
rect 232 -237 233 -236
rect 233 -237 234 -236
rect 234 -237 235 -236
rect 235 -237 236 -236
rect 236 -237 237 -236
rect 237 -237 238 -236
rect 238 -237 239 -236
rect 239 -237 240 -236
rect 240 -237 241 -236
rect 241 -237 242 -236
rect 242 -237 243 -236
rect 243 -237 244 -236
rect 244 -237 245 -236
rect 245 -237 246 -236
rect 246 -237 247 -236
rect 247 -237 248 -236
rect 248 -237 249 -236
rect 249 -237 250 -236
rect 250 -237 251 -236
rect 251 -237 252 -236
rect 252 -237 253 -236
rect 253 -237 254 -236
rect 254 -237 255 -236
rect 255 -237 256 -236
rect 256 -237 257 -236
rect 257 -237 258 -236
rect 258 -237 259 -236
rect 259 -237 260 -236
rect 260 -237 261 -236
rect 261 -237 262 -236
rect 262 -237 263 -236
rect 263 -237 264 -236
rect 264 -237 265 -236
rect 265 -237 266 -236
rect 266 -237 267 -236
rect 267 -237 268 -236
rect 268 -237 269 -236
rect 269 -237 270 -236
rect 270 -237 271 -236
rect 271 -237 272 -236
rect 272 -237 273 -236
rect 273 -237 274 -236
rect 274 -237 275 -236
rect 275 -237 276 -236
rect 276 -237 277 -236
rect 277 -237 278 -236
rect 278 -237 279 -236
rect 279 -237 280 -236
rect 280 -237 281 -236
rect 281 -237 282 -236
rect 282 -237 283 -236
rect 283 -237 284 -236
rect 284 -237 285 -236
rect 285 -237 286 -236
rect 286 -237 287 -236
rect 287 -237 288 -236
rect 288 -237 289 -236
rect 289 -237 290 -236
rect 290 -237 291 -236
rect 291 -237 292 -236
rect 292 -237 293 -236
rect 293 -237 294 -236
rect 294 -237 295 -236
rect 295 -237 296 -236
rect 296 -237 297 -236
rect 297 -237 298 -236
rect 298 -237 299 -236
rect 299 -237 300 -236
rect 300 -237 301 -236
rect 301 -237 302 -236
rect 302 -237 303 -236
rect 303 -237 304 -236
rect 304 -237 305 -236
rect 305 -237 306 -236
rect 306 -237 307 -236
rect 307 -237 308 -236
rect 308 -237 309 -236
rect 309 -237 310 -236
rect 310 -237 311 -236
rect 311 -237 312 -236
rect 312 -237 313 -236
rect 313 -237 314 -236
rect 314 -237 315 -236
rect 315 -237 316 -236
rect 316 -237 317 -236
rect 317 -237 318 -236
rect 318 -237 319 -236
rect 319 -237 320 -236
rect 320 -237 321 -236
rect 321 -237 322 -236
rect 322 -237 323 -236
rect 323 -237 324 -236
rect 324 -237 325 -236
rect 325 -237 326 -236
rect 326 -237 327 -236
rect 327 -237 328 -236
rect 328 -237 329 -236
rect 329 -237 330 -236
rect 330 -237 331 -236
rect 331 -237 332 -236
rect 332 -237 333 -236
rect 333 -237 334 -236
rect 334 -237 335 -236
rect 335 -237 336 -236
rect 336 -237 337 -236
rect 337 -237 338 -236
rect 338 -237 339 -236
rect 339 -237 340 -236
rect 340 -237 341 -236
rect 341 -237 342 -236
rect 342 -237 343 -236
rect 343 -237 344 -236
rect 344 -237 345 -236
rect 345 -237 346 -236
rect 346 -237 347 -236
rect 347 -237 348 -236
rect 348 -237 349 -236
rect 349 -237 350 -236
rect 350 -237 351 -236
rect 351 -237 352 -236
rect 352 -237 353 -236
rect 353 -237 354 -236
rect 354 -237 355 -236
rect 355 -237 356 -236
rect 356 -237 357 -236
rect 357 -237 358 -236
rect 358 -237 359 -236
rect 359 -237 360 -236
rect 360 -237 361 -236
rect 361 -237 362 -236
rect 362 -237 363 -236
rect 363 -237 364 -236
rect 364 -237 365 -236
rect 365 -237 366 -236
rect 366 -237 367 -236
rect 367 -237 368 -236
rect 368 -237 369 -236
rect 369 -237 370 -236
rect 370 -237 371 -236
rect 371 -237 372 -236
rect 372 -237 373 -236
rect 373 -237 374 -236
rect 374 -237 375 -236
rect 375 -237 376 -236
rect 376 -237 377 -236
rect 377 -237 378 -236
rect 378 -237 379 -236
rect 379 -237 380 -236
rect 380 -237 381 -236
rect 381 -237 382 -236
rect 382 -237 383 -236
rect 383 -237 384 -236
rect 384 -237 385 -236
rect 385 -237 386 -236
rect 386 -237 387 -236
rect 387 -237 388 -236
rect 388 -237 389 -236
rect 389 -237 390 -236
rect 390 -237 391 -236
rect 391 -237 392 -236
rect 392 -237 393 -236
rect 393 -237 394 -236
rect 394 -237 395 -236
rect 395 -237 396 -236
rect 396 -237 397 -236
rect 397 -237 398 -236
rect 398 -237 399 -236
rect 399 -237 400 -236
rect 400 -237 401 -236
rect 401 -237 402 -236
rect 402 -237 403 -236
rect 403 -237 404 -236
rect 404 -237 405 -236
rect 405 -237 406 -236
rect 406 -237 407 -236
rect 407 -237 408 -236
rect 408 -237 409 -236
rect 409 -237 410 -236
rect 410 -237 411 -236
rect 411 -237 412 -236
rect 412 -237 413 -236
rect 413 -237 414 -236
rect 414 -237 415 -236
rect 415 -237 416 -236
rect 416 -237 417 -236
rect 417 -237 418 -236
rect 418 -237 419 -236
rect 419 -237 420 -236
rect 420 -237 421 -236
rect 421 -237 422 -236
rect 422 -237 423 -236
rect 423 -237 424 -236
rect 424 -237 425 -236
rect 425 -237 426 -236
rect 426 -237 427 -236
rect 427 -237 428 -236
rect 428 -237 429 -236
rect 429 -237 430 -236
rect 430 -237 431 -236
rect 431 -237 432 -236
rect 432 -237 433 -236
rect 433 -237 434 -236
rect 434 -237 435 -236
rect 435 -237 436 -236
rect 436 -237 437 -236
rect 437 -237 438 -236
rect 438 -237 439 -236
rect 439 -237 440 -236
rect 440 -237 441 -236
rect 441 -237 442 -236
rect 442 -237 443 -236
rect 443 -237 444 -236
rect 444 -237 445 -236
rect 445 -237 446 -236
rect 446 -237 447 -236
rect 447 -237 448 -236
rect 448 -237 449 -236
rect 449 -237 450 -236
rect 450 -237 451 -236
rect 451 -237 452 -236
rect 452 -237 453 -236
rect 453 -237 454 -236
rect 454 -237 455 -236
rect 455 -237 456 -236
rect 456 -237 457 -236
rect 457 -237 458 -236
rect 458 -237 459 -236
rect 459 -237 460 -236
rect 460 -237 461 -236
rect 461 -237 462 -236
rect 462 -237 463 -236
rect 463 -237 464 -236
rect 464 -237 465 -236
rect 465 -237 466 -236
rect 466 -237 467 -236
rect 467 -237 468 -236
rect 468 -237 469 -236
rect 469 -237 470 -236
rect 470 -237 471 -236
rect 471 -237 472 -236
rect 472 -237 473 -236
rect 473 -237 474 -236
rect 474 -237 475 -236
rect 475 -237 476 -236
rect 476 -237 477 -236
rect 477 -237 478 -236
rect 478 -237 479 -236
rect 479 -237 480 -236
rect 2 -238 3 -237
rect 3 -238 4 -237
rect 4 -238 5 -237
rect 5 -238 6 -237
rect 6 -238 7 -237
rect 7 -238 8 -237
rect 8 -238 9 -237
rect 9 -238 10 -237
rect 10 -238 11 -237
rect 11 -238 12 -237
rect 12 -238 13 -237
rect 13 -238 14 -237
rect 14 -238 15 -237
rect 15 -238 16 -237
rect 16 -238 17 -237
rect 17 -238 18 -237
rect 18 -238 19 -237
rect 19 -238 20 -237
rect 20 -238 21 -237
rect 21 -238 22 -237
rect 22 -238 23 -237
rect 23 -238 24 -237
rect 24 -238 25 -237
rect 25 -238 26 -237
rect 26 -238 27 -237
rect 27 -238 28 -237
rect 28 -238 29 -237
rect 29 -238 30 -237
rect 30 -238 31 -237
rect 31 -238 32 -237
rect 32 -238 33 -237
rect 33 -238 34 -237
rect 34 -238 35 -237
rect 35 -238 36 -237
rect 36 -238 37 -237
rect 37 -238 38 -237
rect 38 -238 39 -237
rect 39 -238 40 -237
rect 40 -238 41 -237
rect 41 -238 42 -237
rect 42 -238 43 -237
rect 43 -238 44 -237
rect 44 -238 45 -237
rect 45 -238 46 -237
rect 46 -238 47 -237
rect 47 -238 48 -237
rect 48 -238 49 -237
rect 49 -238 50 -237
rect 50 -238 51 -237
rect 51 -238 52 -237
rect 52 -238 53 -237
rect 53 -238 54 -237
rect 54 -238 55 -237
rect 55 -238 56 -237
rect 56 -238 57 -237
rect 57 -238 58 -237
rect 58 -238 59 -237
rect 59 -238 60 -237
rect 60 -238 61 -237
rect 61 -238 62 -237
rect 62 -238 63 -237
rect 63 -238 64 -237
rect 64 -238 65 -237
rect 65 -238 66 -237
rect 66 -238 67 -237
rect 67 -238 68 -237
rect 68 -238 69 -237
rect 69 -238 70 -237
rect 70 -238 71 -237
rect 71 -238 72 -237
rect 72 -238 73 -237
rect 73 -238 74 -237
rect 74 -238 75 -237
rect 75 -238 76 -237
rect 76 -238 77 -237
rect 77 -238 78 -237
rect 78 -238 79 -237
rect 79 -238 80 -237
rect 80 -238 81 -237
rect 81 -238 82 -237
rect 82 -238 83 -237
rect 83 -238 84 -237
rect 84 -238 85 -237
rect 85 -238 86 -237
rect 86 -238 87 -237
rect 87 -238 88 -237
rect 88 -238 89 -237
rect 89 -238 90 -237
rect 90 -238 91 -237
rect 91 -238 92 -237
rect 92 -238 93 -237
rect 93 -238 94 -237
rect 94 -238 95 -237
rect 95 -238 96 -237
rect 96 -238 97 -237
rect 97 -238 98 -237
rect 98 -238 99 -237
rect 99 -238 100 -237
rect 100 -238 101 -237
rect 101 -238 102 -237
rect 102 -238 103 -237
rect 103 -238 104 -237
rect 104 -238 105 -237
rect 105 -238 106 -237
rect 106 -238 107 -237
rect 107 -238 108 -237
rect 108 -238 109 -237
rect 109 -238 110 -237
rect 110 -238 111 -237
rect 111 -238 112 -237
rect 112 -238 113 -237
rect 113 -238 114 -237
rect 114 -238 115 -237
rect 115 -238 116 -237
rect 116 -238 117 -237
rect 117 -238 118 -237
rect 118 -238 119 -237
rect 119 -238 120 -237
rect 120 -238 121 -237
rect 121 -238 122 -237
rect 122 -238 123 -237
rect 123 -238 124 -237
rect 124 -238 125 -237
rect 125 -238 126 -237
rect 126 -238 127 -237
rect 127 -238 128 -237
rect 128 -238 129 -237
rect 129 -238 130 -237
rect 130 -238 131 -237
rect 131 -238 132 -237
rect 132 -238 133 -237
rect 133 -238 134 -237
rect 134 -238 135 -237
rect 135 -238 136 -237
rect 136 -238 137 -237
rect 137 -238 138 -237
rect 138 -238 139 -237
rect 139 -238 140 -237
rect 140 -238 141 -237
rect 141 -238 142 -237
rect 142 -238 143 -237
rect 143 -238 144 -237
rect 144 -238 145 -237
rect 145 -238 146 -237
rect 146 -238 147 -237
rect 147 -238 148 -237
rect 148 -238 149 -237
rect 149 -238 150 -237
rect 150 -238 151 -237
rect 151 -238 152 -237
rect 152 -238 153 -237
rect 153 -238 154 -237
rect 154 -238 155 -237
rect 155 -238 156 -237
rect 156 -238 157 -237
rect 157 -238 158 -237
rect 158 -238 159 -237
rect 159 -238 160 -237
rect 160 -238 161 -237
rect 161 -238 162 -237
rect 162 -238 163 -237
rect 163 -238 164 -237
rect 164 -238 165 -237
rect 165 -238 166 -237
rect 166 -238 167 -237
rect 167 -238 168 -237
rect 168 -238 169 -237
rect 169 -238 170 -237
rect 170 -238 171 -237
rect 171 -238 172 -237
rect 172 -238 173 -237
rect 173 -238 174 -237
rect 174 -238 175 -237
rect 175 -238 176 -237
rect 176 -238 177 -237
rect 177 -238 178 -237
rect 178 -238 179 -237
rect 179 -238 180 -237
rect 180 -238 181 -237
rect 181 -238 182 -237
rect 182 -238 183 -237
rect 183 -238 184 -237
rect 184 -238 185 -237
rect 185 -238 186 -237
rect 186 -238 187 -237
rect 187 -238 188 -237
rect 188 -238 189 -237
rect 189 -238 190 -237
rect 190 -238 191 -237
rect 191 -238 192 -237
rect 192 -238 193 -237
rect 193 -238 194 -237
rect 194 -238 195 -237
rect 195 -238 196 -237
rect 196 -238 197 -237
rect 197 -238 198 -237
rect 198 -238 199 -237
rect 199 -238 200 -237
rect 200 -238 201 -237
rect 201 -238 202 -237
rect 202 -238 203 -237
rect 203 -238 204 -237
rect 204 -238 205 -237
rect 205 -238 206 -237
rect 206 -238 207 -237
rect 207 -238 208 -237
rect 208 -238 209 -237
rect 209 -238 210 -237
rect 210 -238 211 -237
rect 211 -238 212 -237
rect 212 -238 213 -237
rect 213 -238 214 -237
rect 214 -238 215 -237
rect 215 -238 216 -237
rect 216 -238 217 -237
rect 217 -238 218 -237
rect 218 -238 219 -237
rect 219 -238 220 -237
rect 220 -238 221 -237
rect 221 -238 222 -237
rect 222 -238 223 -237
rect 223 -238 224 -237
rect 224 -238 225 -237
rect 225 -238 226 -237
rect 226 -238 227 -237
rect 227 -238 228 -237
rect 228 -238 229 -237
rect 229 -238 230 -237
rect 230 -238 231 -237
rect 231 -238 232 -237
rect 232 -238 233 -237
rect 233 -238 234 -237
rect 234 -238 235 -237
rect 235 -238 236 -237
rect 236 -238 237 -237
rect 237 -238 238 -237
rect 238 -238 239 -237
rect 239 -238 240 -237
rect 240 -238 241 -237
rect 241 -238 242 -237
rect 242 -238 243 -237
rect 243 -238 244 -237
rect 244 -238 245 -237
rect 245 -238 246 -237
rect 246 -238 247 -237
rect 247 -238 248 -237
rect 248 -238 249 -237
rect 249 -238 250 -237
rect 250 -238 251 -237
rect 251 -238 252 -237
rect 252 -238 253 -237
rect 253 -238 254 -237
rect 254 -238 255 -237
rect 255 -238 256 -237
rect 256 -238 257 -237
rect 257 -238 258 -237
rect 258 -238 259 -237
rect 259 -238 260 -237
rect 260 -238 261 -237
rect 261 -238 262 -237
rect 262 -238 263 -237
rect 263 -238 264 -237
rect 264 -238 265 -237
rect 265 -238 266 -237
rect 266 -238 267 -237
rect 267 -238 268 -237
rect 268 -238 269 -237
rect 269 -238 270 -237
rect 270 -238 271 -237
rect 271 -238 272 -237
rect 272 -238 273 -237
rect 273 -238 274 -237
rect 274 -238 275 -237
rect 275 -238 276 -237
rect 276 -238 277 -237
rect 277 -238 278 -237
rect 278 -238 279 -237
rect 279 -238 280 -237
rect 280 -238 281 -237
rect 281 -238 282 -237
rect 282 -238 283 -237
rect 283 -238 284 -237
rect 284 -238 285 -237
rect 285 -238 286 -237
rect 286 -238 287 -237
rect 287 -238 288 -237
rect 288 -238 289 -237
rect 289 -238 290 -237
rect 290 -238 291 -237
rect 291 -238 292 -237
rect 292 -238 293 -237
rect 293 -238 294 -237
rect 294 -238 295 -237
rect 295 -238 296 -237
rect 296 -238 297 -237
rect 297 -238 298 -237
rect 298 -238 299 -237
rect 299 -238 300 -237
rect 300 -238 301 -237
rect 301 -238 302 -237
rect 302 -238 303 -237
rect 303 -238 304 -237
rect 304 -238 305 -237
rect 305 -238 306 -237
rect 306 -238 307 -237
rect 307 -238 308 -237
rect 308 -238 309 -237
rect 309 -238 310 -237
rect 310 -238 311 -237
rect 311 -238 312 -237
rect 312 -238 313 -237
rect 313 -238 314 -237
rect 314 -238 315 -237
rect 315 -238 316 -237
rect 316 -238 317 -237
rect 317 -238 318 -237
rect 318 -238 319 -237
rect 319 -238 320 -237
rect 320 -238 321 -237
rect 321 -238 322 -237
rect 322 -238 323 -237
rect 323 -238 324 -237
rect 324 -238 325 -237
rect 325 -238 326 -237
rect 326 -238 327 -237
rect 327 -238 328 -237
rect 328 -238 329 -237
rect 329 -238 330 -237
rect 330 -238 331 -237
rect 331 -238 332 -237
rect 332 -238 333 -237
rect 333 -238 334 -237
rect 334 -238 335 -237
rect 335 -238 336 -237
rect 336 -238 337 -237
rect 337 -238 338 -237
rect 338 -238 339 -237
rect 339 -238 340 -237
rect 340 -238 341 -237
rect 341 -238 342 -237
rect 342 -238 343 -237
rect 343 -238 344 -237
rect 344 -238 345 -237
rect 345 -238 346 -237
rect 346 -238 347 -237
rect 347 -238 348 -237
rect 348 -238 349 -237
rect 349 -238 350 -237
rect 350 -238 351 -237
rect 351 -238 352 -237
rect 352 -238 353 -237
rect 353 -238 354 -237
rect 354 -238 355 -237
rect 355 -238 356 -237
rect 356 -238 357 -237
rect 357 -238 358 -237
rect 358 -238 359 -237
rect 359 -238 360 -237
rect 360 -238 361 -237
rect 361 -238 362 -237
rect 362 -238 363 -237
rect 363 -238 364 -237
rect 364 -238 365 -237
rect 365 -238 366 -237
rect 366 -238 367 -237
rect 367 -238 368 -237
rect 368 -238 369 -237
rect 369 -238 370 -237
rect 370 -238 371 -237
rect 371 -238 372 -237
rect 372 -238 373 -237
rect 373 -238 374 -237
rect 374 -238 375 -237
rect 375 -238 376 -237
rect 376 -238 377 -237
rect 377 -238 378 -237
rect 378 -238 379 -237
rect 379 -238 380 -237
rect 380 -238 381 -237
rect 381 -238 382 -237
rect 382 -238 383 -237
rect 383 -238 384 -237
rect 384 -238 385 -237
rect 385 -238 386 -237
rect 386 -238 387 -237
rect 387 -238 388 -237
rect 388 -238 389 -237
rect 389 -238 390 -237
rect 390 -238 391 -237
rect 391 -238 392 -237
rect 392 -238 393 -237
rect 393 -238 394 -237
rect 394 -238 395 -237
rect 395 -238 396 -237
rect 396 -238 397 -237
rect 397 -238 398 -237
rect 398 -238 399 -237
rect 399 -238 400 -237
rect 400 -238 401 -237
rect 401 -238 402 -237
rect 402 -238 403 -237
rect 403 -238 404 -237
rect 404 -238 405 -237
rect 405 -238 406 -237
rect 406 -238 407 -237
rect 407 -238 408 -237
rect 408 -238 409 -237
rect 409 -238 410 -237
rect 410 -238 411 -237
rect 411 -238 412 -237
rect 412 -238 413 -237
rect 413 -238 414 -237
rect 414 -238 415 -237
rect 415 -238 416 -237
rect 416 -238 417 -237
rect 417 -238 418 -237
rect 418 -238 419 -237
rect 419 -238 420 -237
rect 420 -238 421 -237
rect 421 -238 422 -237
rect 422 -238 423 -237
rect 423 -238 424 -237
rect 424 -238 425 -237
rect 425 -238 426 -237
rect 426 -238 427 -237
rect 427 -238 428 -237
rect 428 -238 429 -237
rect 429 -238 430 -237
rect 430 -238 431 -237
rect 431 -238 432 -237
rect 432 -238 433 -237
rect 433 -238 434 -237
rect 434 -238 435 -237
rect 435 -238 436 -237
rect 436 -238 437 -237
rect 437 -238 438 -237
rect 438 -238 439 -237
rect 439 -238 440 -237
rect 440 -238 441 -237
rect 441 -238 442 -237
rect 442 -238 443 -237
rect 443 -238 444 -237
rect 444 -238 445 -237
rect 445 -238 446 -237
rect 446 -238 447 -237
rect 447 -238 448 -237
rect 448 -238 449 -237
rect 449 -238 450 -237
rect 450 -238 451 -237
rect 451 -238 452 -237
rect 452 -238 453 -237
rect 453 -238 454 -237
rect 454 -238 455 -237
rect 455 -238 456 -237
rect 456 -238 457 -237
rect 457 -238 458 -237
rect 458 -238 459 -237
rect 459 -238 460 -237
rect 460 -238 461 -237
rect 461 -238 462 -237
rect 462 -238 463 -237
rect 463 -238 464 -237
rect 464 -238 465 -237
rect 465 -238 466 -237
rect 466 -238 467 -237
rect 467 -238 468 -237
rect 468 -238 469 -237
rect 469 -238 470 -237
rect 470 -238 471 -237
rect 471 -238 472 -237
rect 472 -238 473 -237
rect 473 -238 474 -237
rect 474 -238 475 -237
rect 475 -238 476 -237
rect 476 -238 477 -237
rect 477 -238 478 -237
rect 478 -238 479 -237
rect 479 -238 480 -237
rect 2 -239 3 -238
rect 3 -239 4 -238
rect 4 -239 5 -238
rect 5 -239 6 -238
rect 6 -239 7 -238
rect 7 -239 8 -238
rect 8 -239 9 -238
rect 9 -239 10 -238
rect 10 -239 11 -238
rect 11 -239 12 -238
rect 12 -239 13 -238
rect 13 -239 14 -238
rect 14 -239 15 -238
rect 15 -239 16 -238
rect 16 -239 17 -238
rect 17 -239 18 -238
rect 18 -239 19 -238
rect 19 -239 20 -238
rect 20 -239 21 -238
rect 21 -239 22 -238
rect 22 -239 23 -238
rect 23 -239 24 -238
rect 24 -239 25 -238
rect 25 -239 26 -238
rect 26 -239 27 -238
rect 27 -239 28 -238
rect 28 -239 29 -238
rect 29 -239 30 -238
rect 30 -239 31 -238
rect 31 -239 32 -238
rect 32 -239 33 -238
rect 33 -239 34 -238
rect 34 -239 35 -238
rect 35 -239 36 -238
rect 36 -239 37 -238
rect 37 -239 38 -238
rect 38 -239 39 -238
rect 39 -239 40 -238
rect 40 -239 41 -238
rect 41 -239 42 -238
rect 42 -239 43 -238
rect 43 -239 44 -238
rect 44 -239 45 -238
rect 45 -239 46 -238
rect 46 -239 47 -238
rect 47 -239 48 -238
rect 48 -239 49 -238
rect 49 -239 50 -238
rect 50 -239 51 -238
rect 51 -239 52 -238
rect 52 -239 53 -238
rect 53 -239 54 -238
rect 54 -239 55 -238
rect 55 -239 56 -238
rect 56 -239 57 -238
rect 57 -239 58 -238
rect 58 -239 59 -238
rect 59 -239 60 -238
rect 60 -239 61 -238
rect 61 -239 62 -238
rect 62 -239 63 -238
rect 63 -239 64 -238
rect 64 -239 65 -238
rect 65 -239 66 -238
rect 66 -239 67 -238
rect 67 -239 68 -238
rect 68 -239 69 -238
rect 69 -239 70 -238
rect 70 -239 71 -238
rect 71 -239 72 -238
rect 72 -239 73 -238
rect 73 -239 74 -238
rect 74 -239 75 -238
rect 75 -239 76 -238
rect 76 -239 77 -238
rect 77 -239 78 -238
rect 78 -239 79 -238
rect 79 -239 80 -238
rect 80 -239 81 -238
rect 81 -239 82 -238
rect 82 -239 83 -238
rect 83 -239 84 -238
rect 84 -239 85 -238
rect 85 -239 86 -238
rect 86 -239 87 -238
rect 87 -239 88 -238
rect 88 -239 89 -238
rect 89 -239 90 -238
rect 90 -239 91 -238
rect 91 -239 92 -238
rect 92 -239 93 -238
rect 93 -239 94 -238
rect 94 -239 95 -238
rect 95 -239 96 -238
rect 96 -239 97 -238
rect 97 -239 98 -238
rect 98 -239 99 -238
rect 99 -239 100 -238
rect 100 -239 101 -238
rect 101 -239 102 -238
rect 102 -239 103 -238
rect 103 -239 104 -238
rect 104 -239 105 -238
rect 105 -239 106 -238
rect 106 -239 107 -238
rect 107 -239 108 -238
rect 108 -239 109 -238
rect 109 -239 110 -238
rect 110 -239 111 -238
rect 111 -239 112 -238
rect 112 -239 113 -238
rect 113 -239 114 -238
rect 114 -239 115 -238
rect 115 -239 116 -238
rect 116 -239 117 -238
rect 117 -239 118 -238
rect 118 -239 119 -238
rect 119 -239 120 -238
rect 120 -239 121 -238
rect 121 -239 122 -238
rect 122 -239 123 -238
rect 123 -239 124 -238
rect 124 -239 125 -238
rect 125 -239 126 -238
rect 126 -239 127 -238
rect 127 -239 128 -238
rect 128 -239 129 -238
rect 129 -239 130 -238
rect 130 -239 131 -238
rect 131 -239 132 -238
rect 132 -239 133 -238
rect 133 -239 134 -238
rect 134 -239 135 -238
rect 135 -239 136 -238
rect 136 -239 137 -238
rect 137 -239 138 -238
rect 138 -239 139 -238
rect 139 -239 140 -238
rect 140 -239 141 -238
rect 141 -239 142 -238
rect 142 -239 143 -238
rect 143 -239 144 -238
rect 144 -239 145 -238
rect 145 -239 146 -238
rect 146 -239 147 -238
rect 147 -239 148 -238
rect 148 -239 149 -238
rect 149 -239 150 -238
rect 150 -239 151 -238
rect 151 -239 152 -238
rect 152 -239 153 -238
rect 153 -239 154 -238
rect 154 -239 155 -238
rect 155 -239 156 -238
rect 156 -239 157 -238
rect 157 -239 158 -238
rect 158 -239 159 -238
rect 159 -239 160 -238
rect 160 -239 161 -238
rect 161 -239 162 -238
rect 162 -239 163 -238
rect 163 -239 164 -238
rect 164 -239 165 -238
rect 165 -239 166 -238
rect 166 -239 167 -238
rect 167 -239 168 -238
rect 168 -239 169 -238
rect 169 -239 170 -238
rect 170 -239 171 -238
rect 171 -239 172 -238
rect 172 -239 173 -238
rect 173 -239 174 -238
rect 174 -239 175 -238
rect 175 -239 176 -238
rect 176 -239 177 -238
rect 177 -239 178 -238
rect 178 -239 179 -238
rect 179 -239 180 -238
rect 180 -239 181 -238
rect 181 -239 182 -238
rect 182 -239 183 -238
rect 183 -239 184 -238
rect 184 -239 185 -238
rect 185 -239 186 -238
rect 186 -239 187 -238
rect 187 -239 188 -238
rect 188 -239 189 -238
rect 189 -239 190 -238
rect 190 -239 191 -238
rect 191 -239 192 -238
rect 192 -239 193 -238
rect 193 -239 194 -238
rect 194 -239 195 -238
rect 195 -239 196 -238
rect 196 -239 197 -238
rect 197 -239 198 -238
rect 198 -239 199 -238
rect 199 -239 200 -238
rect 200 -239 201 -238
rect 201 -239 202 -238
rect 202 -239 203 -238
rect 203 -239 204 -238
rect 204 -239 205 -238
rect 205 -239 206 -238
rect 206 -239 207 -238
rect 207 -239 208 -238
rect 208 -239 209 -238
rect 209 -239 210 -238
rect 210 -239 211 -238
rect 211 -239 212 -238
rect 212 -239 213 -238
rect 213 -239 214 -238
rect 214 -239 215 -238
rect 215 -239 216 -238
rect 216 -239 217 -238
rect 217 -239 218 -238
rect 218 -239 219 -238
rect 219 -239 220 -238
rect 220 -239 221 -238
rect 221 -239 222 -238
rect 222 -239 223 -238
rect 223 -239 224 -238
rect 224 -239 225 -238
rect 225 -239 226 -238
rect 226 -239 227 -238
rect 227 -239 228 -238
rect 228 -239 229 -238
rect 229 -239 230 -238
rect 230 -239 231 -238
rect 231 -239 232 -238
rect 232 -239 233 -238
rect 233 -239 234 -238
rect 234 -239 235 -238
rect 235 -239 236 -238
rect 236 -239 237 -238
rect 237 -239 238 -238
rect 238 -239 239 -238
rect 239 -239 240 -238
rect 240 -239 241 -238
rect 241 -239 242 -238
rect 242 -239 243 -238
rect 243 -239 244 -238
rect 244 -239 245 -238
rect 245 -239 246 -238
rect 246 -239 247 -238
rect 247 -239 248 -238
rect 248 -239 249 -238
rect 249 -239 250 -238
rect 250 -239 251 -238
rect 251 -239 252 -238
rect 252 -239 253 -238
rect 253 -239 254 -238
rect 254 -239 255 -238
rect 255 -239 256 -238
rect 256 -239 257 -238
rect 257 -239 258 -238
rect 258 -239 259 -238
rect 259 -239 260 -238
rect 260 -239 261 -238
rect 261 -239 262 -238
rect 262 -239 263 -238
rect 263 -239 264 -238
rect 264 -239 265 -238
rect 265 -239 266 -238
rect 266 -239 267 -238
rect 267 -239 268 -238
rect 268 -239 269 -238
rect 269 -239 270 -238
rect 270 -239 271 -238
rect 271 -239 272 -238
rect 272 -239 273 -238
rect 273 -239 274 -238
rect 274 -239 275 -238
rect 275 -239 276 -238
rect 276 -239 277 -238
rect 277 -239 278 -238
rect 278 -239 279 -238
rect 279 -239 280 -238
rect 280 -239 281 -238
rect 281 -239 282 -238
rect 282 -239 283 -238
rect 283 -239 284 -238
rect 284 -239 285 -238
rect 285 -239 286 -238
rect 286 -239 287 -238
rect 287 -239 288 -238
rect 288 -239 289 -238
rect 289 -239 290 -238
rect 290 -239 291 -238
rect 291 -239 292 -238
rect 292 -239 293 -238
rect 293 -239 294 -238
rect 294 -239 295 -238
rect 295 -239 296 -238
rect 296 -239 297 -238
rect 297 -239 298 -238
rect 298 -239 299 -238
rect 299 -239 300 -238
rect 300 -239 301 -238
rect 301 -239 302 -238
rect 302 -239 303 -238
rect 303 -239 304 -238
rect 304 -239 305 -238
rect 305 -239 306 -238
rect 306 -239 307 -238
rect 307 -239 308 -238
rect 308 -239 309 -238
rect 309 -239 310 -238
rect 310 -239 311 -238
rect 311 -239 312 -238
rect 312 -239 313 -238
rect 313 -239 314 -238
rect 314 -239 315 -238
rect 315 -239 316 -238
rect 316 -239 317 -238
rect 317 -239 318 -238
rect 318 -239 319 -238
rect 319 -239 320 -238
rect 320 -239 321 -238
rect 321 -239 322 -238
rect 322 -239 323 -238
rect 323 -239 324 -238
rect 324 -239 325 -238
rect 325 -239 326 -238
rect 326 -239 327 -238
rect 327 -239 328 -238
rect 328 -239 329 -238
rect 329 -239 330 -238
rect 330 -239 331 -238
rect 331 -239 332 -238
rect 332 -239 333 -238
rect 333 -239 334 -238
rect 334 -239 335 -238
rect 335 -239 336 -238
rect 336 -239 337 -238
rect 337 -239 338 -238
rect 338 -239 339 -238
rect 339 -239 340 -238
rect 340 -239 341 -238
rect 341 -239 342 -238
rect 342 -239 343 -238
rect 343 -239 344 -238
rect 344 -239 345 -238
rect 345 -239 346 -238
rect 346 -239 347 -238
rect 347 -239 348 -238
rect 348 -239 349 -238
rect 349 -239 350 -238
rect 350 -239 351 -238
rect 351 -239 352 -238
rect 352 -239 353 -238
rect 353 -239 354 -238
rect 354 -239 355 -238
rect 355 -239 356 -238
rect 356 -239 357 -238
rect 357 -239 358 -238
rect 358 -239 359 -238
rect 359 -239 360 -238
rect 360 -239 361 -238
rect 361 -239 362 -238
rect 362 -239 363 -238
rect 363 -239 364 -238
rect 364 -239 365 -238
rect 365 -239 366 -238
rect 366 -239 367 -238
rect 367 -239 368 -238
rect 368 -239 369 -238
rect 369 -239 370 -238
rect 370 -239 371 -238
rect 371 -239 372 -238
rect 372 -239 373 -238
rect 373 -239 374 -238
rect 374 -239 375 -238
rect 375 -239 376 -238
rect 376 -239 377 -238
rect 377 -239 378 -238
rect 378 -239 379 -238
rect 379 -239 380 -238
rect 380 -239 381 -238
rect 381 -239 382 -238
rect 382 -239 383 -238
rect 383 -239 384 -238
rect 384 -239 385 -238
rect 385 -239 386 -238
rect 386 -239 387 -238
rect 387 -239 388 -238
rect 388 -239 389 -238
rect 389 -239 390 -238
rect 390 -239 391 -238
rect 391 -239 392 -238
rect 392 -239 393 -238
rect 393 -239 394 -238
rect 394 -239 395 -238
rect 395 -239 396 -238
rect 396 -239 397 -238
rect 397 -239 398 -238
rect 398 -239 399 -238
rect 399 -239 400 -238
rect 400 -239 401 -238
rect 401 -239 402 -238
rect 402 -239 403 -238
rect 403 -239 404 -238
rect 404 -239 405 -238
rect 405 -239 406 -238
rect 406 -239 407 -238
rect 407 -239 408 -238
rect 408 -239 409 -238
rect 409 -239 410 -238
rect 410 -239 411 -238
rect 411 -239 412 -238
rect 412 -239 413 -238
rect 413 -239 414 -238
rect 414 -239 415 -238
rect 415 -239 416 -238
rect 416 -239 417 -238
rect 417 -239 418 -238
rect 418 -239 419 -238
rect 419 -239 420 -238
rect 420 -239 421 -238
rect 421 -239 422 -238
rect 422 -239 423 -238
rect 423 -239 424 -238
rect 424 -239 425 -238
rect 425 -239 426 -238
rect 426 -239 427 -238
rect 427 -239 428 -238
rect 428 -239 429 -238
rect 429 -239 430 -238
rect 430 -239 431 -238
rect 431 -239 432 -238
rect 432 -239 433 -238
rect 433 -239 434 -238
rect 434 -239 435 -238
rect 435 -239 436 -238
rect 436 -239 437 -238
rect 437 -239 438 -238
rect 438 -239 439 -238
rect 439 -239 440 -238
rect 440 -239 441 -238
rect 441 -239 442 -238
rect 442 -239 443 -238
rect 443 -239 444 -238
rect 444 -239 445 -238
rect 445 -239 446 -238
rect 446 -239 447 -238
rect 447 -239 448 -238
rect 448 -239 449 -238
rect 449 -239 450 -238
rect 450 -239 451 -238
rect 451 -239 452 -238
rect 452 -239 453 -238
rect 453 -239 454 -238
rect 454 -239 455 -238
rect 455 -239 456 -238
rect 456 -239 457 -238
rect 457 -239 458 -238
rect 458 -239 459 -238
rect 459 -239 460 -238
rect 460 -239 461 -238
rect 461 -239 462 -238
rect 462 -239 463 -238
rect 463 -239 464 -238
rect 464 -239 465 -238
rect 465 -239 466 -238
rect 466 -239 467 -238
rect 467 -239 468 -238
rect 468 -239 469 -238
rect 469 -239 470 -238
rect 470 -239 471 -238
rect 471 -239 472 -238
rect 472 -239 473 -238
rect 473 -239 474 -238
rect 474 -239 475 -238
rect 475 -239 476 -238
rect 476 -239 477 -238
rect 477 -239 478 -238
rect 478 -239 479 -238
rect 479 -239 480 -238
rect 2 -240 3 -239
rect 3 -240 4 -239
rect 4 -240 5 -239
rect 5 -240 6 -239
rect 6 -240 7 -239
rect 7 -240 8 -239
rect 8 -240 9 -239
rect 9 -240 10 -239
rect 10 -240 11 -239
rect 11 -240 12 -239
rect 12 -240 13 -239
rect 13 -240 14 -239
rect 14 -240 15 -239
rect 15 -240 16 -239
rect 16 -240 17 -239
rect 17 -240 18 -239
rect 18 -240 19 -239
rect 19 -240 20 -239
rect 20 -240 21 -239
rect 21 -240 22 -239
rect 22 -240 23 -239
rect 23 -240 24 -239
rect 24 -240 25 -239
rect 25 -240 26 -239
rect 26 -240 27 -239
rect 27 -240 28 -239
rect 28 -240 29 -239
rect 29 -240 30 -239
rect 30 -240 31 -239
rect 31 -240 32 -239
rect 32 -240 33 -239
rect 33 -240 34 -239
rect 34 -240 35 -239
rect 35 -240 36 -239
rect 36 -240 37 -239
rect 37 -240 38 -239
rect 38 -240 39 -239
rect 39 -240 40 -239
rect 40 -240 41 -239
rect 41 -240 42 -239
rect 42 -240 43 -239
rect 43 -240 44 -239
rect 44 -240 45 -239
rect 45 -240 46 -239
rect 46 -240 47 -239
rect 47 -240 48 -239
rect 48 -240 49 -239
rect 49 -240 50 -239
rect 50 -240 51 -239
rect 51 -240 52 -239
rect 52 -240 53 -239
rect 53 -240 54 -239
rect 54 -240 55 -239
rect 55 -240 56 -239
rect 56 -240 57 -239
rect 57 -240 58 -239
rect 58 -240 59 -239
rect 59 -240 60 -239
rect 60 -240 61 -239
rect 61 -240 62 -239
rect 62 -240 63 -239
rect 63 -240 64 -239
rect 64 -240 65 -239
rect 65 -240 66 -239
rect 66 -240 67 -239
rect 67 -240 68 -239
rect 68 -240 69 -239
rect 69 -240 70 -239
rect 70 -240 71 -239
rect 71 -240 72 -239
rect 72 -240 73 -239
rect 73 -240 74 -239
rect 74 -240 75 -239
rect 75 -240 76 -239
rect 76 -240 77 -239
rect 77 -240 78 -239
rect 78 -240 79 -239
rect 79 -240 80 -239
rect 80 -240 81 -239
rect 81 -240 82 -239
rect 82 -240 83 -239
rect 83 -240 84 -239
rect 84 -240 85 -239
rect 85 -240 86 -239
rect 86 -240 87 -239
rect 87 -240 88 -239
rect 88 -240 89 -239
rect 89 -240 90 -239
rect 90 -240 91 -239
rect 91 -240 92 -239
rect 92 -240 93 -239
rect 93 -240 94 -239
rect 94 -240 95 -239
rect 95 -240 96 -239
rect 96 -240 97 -239
rect 97 -240 98 -239
rect 98 -240 99 -239
rect 99 -240 100 -239
rect 100 -240 101 -239
rect 101 -240 102 -239
rect 102 -240 103 -239
rect 103 -240 104 -239
rect 104 -240 105 -239
rect 105 -240 106 -239
rect 106 -240 107 -239
rect 107 -240 108 -239
rect 108 -240 109 -239
rect 109 -240 110 -239
rect 110 -240 111 -239
rect 111 -240 112 -239
rect 112 -240 113 -239
rect 113 -240 114 -239
rect 114 -240 115 -239
rect 115 -240 116 -239
rect 116 -240 117 -239
rect 117 -240 118 -239
rect 118 -240 119 -239
rect 119 -240 120 -239
rect 120 -240 121 -239
rect 121 -240 122 -239
rect 122 -240 123 -239
rect 123 -240 124 -239
rect 124 -240 125 -239
rect 125 -240 126 -239
rect 126 -240 127 -239
rect 127 -240 128 -239
rect 128 -240 129 -239
rect 129 -240 130 -239
rect 130 -240 131 -239
rect 131 -240 132 -239
rect 132 -240 133 -239
rect 133 -240 134 -239
rect 134 -240 135 -239
rect 135 -240 136 -239
rect 136 -240 137 -239
rect 137 -240 138 -239
rect 138 -240 139 -239
rect 139 -240 140 -239
rect 140 -240 141 -239
rect 141 -240 142 -239
rect 142 -240 143 -239
rect 143 -240 144 -239
rect 144 -240 145 -239
rect 145 -240 146 -239
rect 146 -240 147 -239
rect 147 -240 148 -239
rect 148 -240 149 -239
rect 149 -240 150 -239
rect 150 -240 151 -239
rect 151 -240 152 -239
rect 152 -240 153 -239
rect 153 -240 154 -239
rect 154 -240 155 -239
rect 155 -240 156 -239
rect 156 -240 157 -239
rect 157 -240 158 -239
rect 158 -240 159 -239
rect 159 -240 160 -239
rect 160 -240 161 -239
rect 161 -240 162 -239
rect 162 -240 163 -239
rect 163 -240 164 -239
rect 164 -240 165 -239
rect 165 -240 166 -239
rect 166 -240 167 -239
rect 167 -240 168 -239
rect 168 -240 169 -239
rect 169 -240 170 -239
rect 170 -240 171 -239
rect 171 -240 172 -239
rect 172 -240 173 -239
rect 173 -240 174 -239
rect 174 -240 175 -239
rect 175 -240 176 -239
rect 176 -240 177 -239
rect 177 -240 178 -239
rect 178 -240 179 -239
rect 179 -240 180 -239
rect 180 -240 181 -239
rect 181 -240 182 -239
rect 182 -240 183 -239
rect 183 -240 184 -239
rect 184 -240 185 -239
rect 185 -240 186 -239
rect 186 -240 187 -239
rect 187 -240 188 -239
rect 188 -240 189 -239
rect 189 -240 190 -239
rect 190 -240 191 -239
rect 191 -240 192 -239
rect 192 -240 193 -239
rect 193 -240 194 -239
rect 194 -240 195 -239
rect 195 -240 196 -239
rect 196 -240 197 -239
rect 197 -240 198 -239
rect 198 -240 199 -239
rect 199 -240 200 -239
rect 200 -240 201 -239
rect 201 -240 202 -239
rect 202 -240 203 -239
rect 203 -240 204 -239
rect 204 -240 205 -239
rect 205 -240 206 -239
rect 206 -240 207 -239
rect 207 -240 208 -239
rect 208 -240 209 -239
rect 209 -240 210 -239
rect 210 -240 211 -239
rect 211 -240 212 -239
rect 212 -240 213 -239
rect 213 -240 214 -239
rect 214 -240 215 -239
rect 215 -240 216 -239
rect 216 -240 217 -239
rect 217 -240 218 -239
rect 218 -240 219 -239
rect 219 -240 220 -239
rect 220 -240 221 -239
rect 221 -240 222 -239
rect 222 -240 223 -239
rect 223 -240 224 -239
rect 224 -240 225 -239
rect 225 -240 226 -239
rect 226 -240 227 -239
rect 227 -240 228 -239
rect 228 -240 229 -239
rect 229 -240 230 -239
rect 230 -240 231 -239
rect 231 -240 232 -239
rect 232 -240 233 -239
rect 233 -240 234 -239
rect 234 -240 235 -239
rect 235 -240 236 -239
rect 236 -240 237 -239
rect 237 -240 238 -239
rect 238 -240 239 -239
rect 239 -240 240 -239
rect 240 -240 241 -239
rect 241 -240 242 -239
rect 242 -240 243 -239
rect 243 -240 244 -239
rect 244 -240 245 -239
rect 245 -240 246 -239
rect 246 -240 247 -239
rect 247 -240 248 -239
rect 248 -240 249 -239
rect 249 -240 250 -239
rect 250 -240 251 -239
rect 251 -240 252 -239
rect 252 -240 253 -239
rect 253 -240 254 -239
rect 254 -240 255 -239
rect 255 -240 256 -239
rect 256 -240 257 -239
rect 257 -240 258 -239
rect 258 -240 259 -239
rect 259 -240 260 -239
rect 260 -240 261 -239
rect 261 -240 262 -239
rect 262 -240 263 -239
rect 263 -240 264 -239
rect 264 -240 265 -239
rect 265 -240 266 -239
rect 266 -240 267 -239
rect 267 -240 268 -239
rect 268 -240 269 -239
rect 269 -240 270 -239
rect 270 -240 271 -239
rect 271 -240 272 -239
rect 272 -240 273 -239
rect 273 -240 274 -239
rect 274 -240 275 -239
rect 275 -240 276 -239
rect 276 -240 277 -239
rect 277 -240 278 -239
rect 278 -240 279 -239
rect 279 -240 280 -239
rect 280 -240 281 -239
rect 281 -240 282 -239
rect 282 -240 283 -239
rect 283 -240 284 -239
rect 284 -240 285 -239
rect 285 -240 286 -239
rect 286 -240 287 -239
rect 287 -240 288 -239
rect 288 -240 289 -239
rect 289 -240 290 -239
rect 290 -240 291 -239
rect 291 -240 292 -239
rect 292 -240 293 -239
rect 293 -240 294 -239
rect 294 -240 295 -239
rect 295 -240 296 -239
rect 296 -240 297 -239
rect 297 -240 298 -239
rect 298 -240 299 -239
rect 299 -240 300 -239
rect 300 -240 301 -239
rect 301 -240 302 -239
rect 302 -240 303 -239
rect 303 -240 304 -239
rect 304 -240 305 -239
rect 305 -240 306 -239
rect 306 -240 307 -239
rect 307 -240 308 -239
rect 308 -240 309 -239
rect 309 -240 310 -239
rect 310 -240 311 -239
rect 311 -240 312 -239
rect 312 -240 313 -239
rect 313 -240 314 -239
rect 314 -240 315 -239
rect 315 -240 316 -239
rect 316 -240 317 -239
rect 317 -240 318 -239
rect 318 -240 319 -239
rect 319 -240 320 -239
rect 320 -240 321 -239
rect 321 -240 322 -239
rect 322 -240 323 -239
rect 323 -240 324 -239
rect 324 -240 325 -239
rect 325 -240 326 -239
rect 326 -240 327 -239
rect 327 -240 328 -239
rect 328 -240 329 -239
rect 329 -240 330 -239
rect 330 -240 331 -239
rect 331 -240 332 -239
rect 332 -240 333 -239
rect 333 -240 334 -239
rect 334 -240 335 -239
rect 335 -240 336 -239
rect 336 -240 337 -239
rect 337 -240 338 -239
rect 338 -240 339 -239
rect 339 -240 340 -239
rect 340 -240 341 -239
rect 341 -240 342 -239
rect 342 -240 343 -239
rect 343 -240 344 -239
rect 344 -240 345 -239
rect 345 -240 346 -239
rect 346 -240 347 -239
rect 347 -240 348 -239
rect 348 -240 349 -239
rect 349 -240 350 -239
rect 350 -240 351 -239
rect 351 -240 352 -239
rect 352 -240 353 -239
rect 353 -240 354 -239
rect 354 -240 355 -239
rect 355 -240 356 -239
rect 356 -240 357 -239
rect 357 -240 358 -239
rect 358 -240 359 -239
rect 359 -240 360 -239
rect 360 -240 361 -239
rect 361 -240 362 -239
rect 362 -240 363 -239
rect 363 -240 364 -239
rect 364 -240 365 -239
rect 365 -240 366 -239
rect 366 -240 367 -239
rect 367 -240 368 -239
rect 368 -240 369 -239
rect 369 -240 370 -239
rect 370 -240 371 -239
rect 371 -240 372 -239
rect 372 -240 373 -239
rect 373 -240 374 -239
rect 374 -240 375 -239
rect 375 -240 376 -239
rect 376 -240 377 -239
rect 377 -240 378 -239
rect 378 -240 379 -239
rect 379 -240 380 -239
rect 380 -240 381 -239
rect 381 -240 382 -239
rect 382 -240 383 -239
rect 383 -240 384 -239
rect 384 -240 385 -239
rect 385 -240 386 -239
rect 386 -240 387 -239
rect 387 -240 388 -239
rect 388 -240 389 -239
rect 389 -240 390 -239
rect 390 -240 391 -239
rect 391 -240 392 -239
rect 392 -240 393 -239
rect 393 -240 394 -239
rect 394 -240 395 -239
rect 395 -240 396 -239
rect 396 -240 397 -239
rect 397 -240 398 -239
rect 398 -240 399 -239
rect 399 -240 400 -239
rect 400 -240 401 -239
rect 401 -240 402 -239
rect 402 -240 403 -239
rect 403 -240 404 -239
rect 404 -240 405 -239
rect 405 -240 406 -239
rect 406 -240 407 -239
rect 407 -240 408 -239
rect 408 -240 409 -239
rect 409 -240 410 -239
rect 410 -240 411 -239
rect 411 -240 412 -239
rect 412 -240 413 -239
rect 413 -240 414 -239
rect 414 -240 415 -239
rect 415 -240 416 -239
rect 416 -240 417 -239
rect 417 -240 418 -239
rect 418 -240 419 -239
rect 419 -240 420 -239
rect 420 -240 421 -239
rect 421 -240 422 -239
rect 422 -240 423 -239
rect 423 -240 424 -239
rect 424 -240 425 -239
rect 425 -240 426 -239
rect 426 -240 427 -239
rect 427 -240 428 -239
rect 428 -240 429 -239
rect 429 -240 430 -239
rect 430 -240 431 -239
rect 431 -240 432 -239
rect 432 -240 433 -239
rect 433 -240 434 -239
rect 434 -240 435 -239
rect 435 -240 436 -239
rect 436 -240 437 -239
rect 437 -240 438 -239
rect 438 -240 439 -239
rect 439 -240 440 -239
rect 440 -240 441 -239
rect 441 -240 442 -239
rect 442 -240 443 -239
rect 443 -240 444 -239
rect 444 -240 445 -239
rect 445 -240 446 -239
rect 446 -240 447 -239
rect 447 -240 448 -239
rect 448 -240 449 -239
rect 449 -240 450 -239
rect 450 -240 451 -239
rect 451 -240 452 -239
rect 452 -240 453 -239
rect 453 -240 454 -239
rect 454 -240 455 -239
rect 455 -240 456 -239
rect 456 -240 457 -239
rect 457 -240 458 -239
rect 458 -240 459 -239
rect 459 -240 460 -239
rect 460 -240 461 -239
rect 461 -240 462 -239
rect 462 -240 463 -239
rect 463 -240 464 -239
rect 464 -240 465 -239
rect 465 -240 466 -239
rect 466 -240 467 -239
rect 467 -240 468 -239
rect 468 -240 469 -239
rect 469 -240 470 -239
rect 470 -240 471 -239
rect 471 -240 472 -239
rect 472 -240 473 -239
rect 473 -240 474 -239
rect 474 -240 475 -239
rect 475 -240 476 -239
rect 476 -240 477 -239
rect 477 -240 478 -239
rect 478 -240 479 -239
rect 479 -240 480 -239
rect 2 -241 3 -240
rect 3 -241 4 -240
rect 4 -241 5 -240
rect 5 -241 6 -240
rect 6 -241 7 -240
rect 7 -241 8 -240
rect 8 -241 9 -240
rect 9 -241 10 -240
rect 10 -241 11 -240
rect 11 -241 12 -240
rect 12 -241 13 -240
rect 13 -241 14 -240
rect 14 -241 15 -240
rect 15 -241 16 -240
rect 16 -241 17 -240
rect 17 -241 18 -240
rect 18 -241 19 -240
rect 19 -241 20 -240
rect 20 -241 21 -240
rect 21 -241 22 -240
rect 22 -241 23 -240
rect 23 -241 24 -240
rect 24 -241 25 -240
rect 25 -241 26 -240
rect 26 -241 27 -240
rect 27 -241 28 -240
rect 28 -241 29 -240
rect 29 -241 30 -240
rect 30 -241 31 -240
rect 31 -241 32 -240
rect 32 -241 33 -240
rect 33 -241 34 -240
rect 34 -241 35 -240
rect 35 -241 36 -240
rect 36 -241 37 -240
rect 37 -241 38 -240
rect 38 -241 39 -240
rect 39 -241 40 -240
rect 40 -241 41 -240
rect 41 -241 42 -240
rect 42 -241 43 -240
rect 43 -241 44 -240
rect 44 -241 45 -240
rect 45 -241 46 -240
rect 46 -241 47 -240
rect 47 -241 48 -240
rect 48 -241 49 -240
rect 49 -241 50 -240
rect 50 -241 51 -240
rect 51 -241 52 -240
rect 52 -241 53 -240
rect 53 -241 54 -240
rect 54 -241 55 -240
rect 55 -241 56 -240
rect 56 -241 57 -240
rect 57 -241 58 -240
rect 58 -241 59 -240
rect 59 -241 60 -240
rect 60 -241 61 -240
rect 61 -241 62 -240
rect 62 -241 63 -240
rect 63 -241 64 -240
rect 64 -241 65 -240
rect 65 -241 66 -240
rect 66 -241 67 -240
rect 67 -241 68 -240
rect 68 -241 69 -240
rect 69 -241 70 -240
rect 70 -241 71 -240
rect 71 -241 72 -240
rect 72 -241 73 -240
rect 73 -241 74 -240
rect 74 -241 75 -240
rect 75 -241 76 -240
rect 76 -241 77 -240
rect 77 -241 78 -240
rect 78 -241 79 -240
rect 79 -241 80 -240
rect 80 -241 81 -240
rect 81 -241 82 -240
rect 82 -241 83 -240
rect 83 -241 84 -240
rect 84 -241 85 -240
rect 85 -241 86 -240
rect 86 -241 87 -240
rect 87 -241 88 -240
rect 88 -241 89 -240
rect 89 -241 90 -240
rect 90 -241 91 -240
rect 91 -241 92 -240
rect 92 -241 93 -240
rect 93 -241 94 -240
rect 94 -241 95 -240
rect 95 -241 96 -240
rect 96 -241 97 -240
rect 97 -241 98 -240
rect 98 -241 99 -240
rect 99 -241 100 -240
rect 100 -241 101 -240
rect 101 -241 102 -240
rect 102 -241 103 -240
rect 103 -241 104 -240
rect 104 -241 105 -240
rect 105 -241 106 -240
rect 106 -241 107 -240
rect 107 -241 108 -240
rect 108 -241 109 -240
rect 109 -241 110 -240
rect 110 -241 111 -240
rect 111 -241 112 -240
rect 112 -241 113 -240
rect 113 -241 114 -240
rect 114 -241 115 -240
rect 115 -241 116 -240
rect 116 -241 117 -240
rect 117 -241 118 -240
rect 118 -241 119 -240
rect 119 -241 120 -240
rect 120 -241 121 -240
rect 121 -241 122 -240
rect 122 -241 123 -240
rect 123 -241 124 -240
rect 124 -241 125 -240
rect 125 -241 126 -240
rect 126 -241 127 -240
rect 127 -241 128 -240
rect 128 -241 129 -240
rect 129 -241 130 -240
rect 130 -241 131 -240
rect 131 -241 132 -240
rect 132 -241 133 -240
rect 133 -241 134 -240
rect 134 -241 135 -240
rect 135 -241 136 -240
rect 136 -241 137 -240
rect 137 -241 138 -240
rect 138 -241 139 -240
rect 139 -241 140 -240
rect 140 -241 141 -240
rect 141 -241 142 -240
rect 142 -241 143 -240
rect 143 -241 144 -240
rect 144 -241 145 -240
rect 145 -241 146 -240
rect 146 -241 147 -240
rect 147 -241 148 -240
rect 148 -241 149 -240
rect 149 -241 150 -240
rect 150 -241 151 -240
rect 151 -241 152 -240
rect 152 -241 153 -240
rect 153 -241 154 -240
rect 154 -241 155 -240
rect 155 -241 156 -240
rect 156 -241 157 -240
rect 157 -241 158 -240
rect 158 -241 159 -240
rect 159 -241 160 -240
rect 160 -241 161 -240
rect 161 -241 162 -240
rect 162 -241 163 -240
rect 163 -241 164 -240
rect 164 -241 165 -240
rect 165 -241 166 -240
rect 166 -241 167 -240
rect 167 -241 168 -240
rect 168 -241 169 -240
rect 169 -241 170 -240
rect 170 -241 171 -240
rect 171 -241 172 -240
rect 172 -241 173 -240
rect 173 -241 174 -240
rect 174 -241 175 -240
rect 175 -241 176 -240
rect 176 -241 177 -240
rect 177 -241 178 -240
rect 178 -241 179 -240
rect 179 -241 180 -240
rect 180 -241 181 -240
rect 181 -241 182 -240
rect 182 -241 183 -240
rect 183 -241 184 -240
rect 184 -241 185 -240
rect 185 -241 186 -240
rect 186 -241 187 -240
rect 187 -241 188 -240
rect 188 -241 189 -240
rect 189 -241 190 -240
rect 190 -241 191 -240
rect 191 -241 192 -240
rect 192 -241 193 -240
rect 193 -241 194 -240
rect 194 -241 195 -240
rect 195 -241 196 -240
rect 196 -241 197 -240
rect 197 -241 198 -240
rect 198 -241 199 -240
rect 199 -241 200 -240
rect 200 -241 201 -240
rect 201 -241 202 -240
rect 202 -241 203 -240
rect 203 -241 204 -240
rect 204 -241 205 -240
rect 205 -241 206 -240
rect 206 -241 207 -240
rect 207 -241 208 -240
rect 208 -241 209 -240
rect 209 -241 210 -240
rect 210 -241 211 -240
rect 211 -241 212 -240
rect 212 -241 213 -240
rect 213 -241 214 -240
rect 214 -241 215 -240
rect 215 -241 216 -240
rect 216 -241 217 -240
rect 217 -241 218 -240
rect 218 -241 219 -240
rect 219 -241 220 -240
rect 220 -241 221 -240
rect 221 -241 222 -240
rect 222 -241 223 -240
rect 223 -241 224 -240
rect 224 -241 225 -240
rect 225 -241 226 -240
rect 226 -241 227 -240
rect 227 -241 228 -240
rect 228 -241 229 -240
rect 229 -241 230 -240
rect 230 -241 231 -240
rect 231 -241 232 -240
rect 232 -241 233 -240
rect 233 -241 234 -240
rect 234 -241 235 -240
rect 235 -241 236 -240
rect 236 -241 237 -240
rect 237 -241 238 -240
rect 238 -241 239 -240
rect 239 -241 240 -240
rect 240 -241 241 -240
rect 241 -241 242 -240
rect 242 -241 243 -240
rect 243 -241 244 -240
rect 244 -241 245 -240
rect 245 -241 246 -240
rect 246 -241 247 -240
rect 247 -241 248 -240
rect 248 -241 249 -240
rect 249 -241 250 -240
rect 250 -241 251 -240
rect 251 -241 252 -240
rect 252 -241 253 -240
rect 253 -241 254 -240
rect 254 -241 255 -240
rect 255 -241 256 -240
rect 256 -241 257 -240
rect 257 -241 258 -240
rect 258 -241 259 -240
rect 259 -241 260 -240
rect 260 -241 261 -240
rect 261 -241 262 -240
rect 262 -241 263 -240
rect 263 -241 264 -240
rect 264 -241 265 -240
rect 265 -241 266 -240
rect 266 -241 267 -240
rect 267 -241 268 -240
rect 268 -241 269 -240
rect 269 -241 270 -240
rect 270 -241 271 -240
rect 271 -241 272 -240
rect 272 -241 273 -240
rect 273 -241 274 -240
rect 274 -241 275 -240
rect 275 -241 276 -240
rect 276 -241 277 -240
rect 277 -241 278 -240
rect 278 -241 279 -240
rect 279 -241 280 -240
rect 280 -241 281 -240
rect 281 -241 282 -240
rect 282 -241 283 -240
rect 283 -241 284 -240
rect 284 -241 285 -240
rect 285 -241 286 -240
rect 286 -241 287 -240
rect 287 -241 288 -240
rect 288 -241 289 -240
rect 289 -241 290 -240
rect 290 -241 291 -240
rect 291 -241 292 -240
rect 292 -241 293 -240
rect 293 -241 294 -240
rect 294 -241 295 -240
rect 295 -241 296 -240
rect 296 -241 297 -240
rect 297 -241 298 -240
rect 298 -241 299 -240
rect 299 -241 300 -240
rect 300 -241 301 -240
rect 301 -241 302 -240
rect 302 -241 303 -240
rect 303 -241 304 -240
rect 304 -241 305 -240
rect 305 -241 306 -240
rect 306 -241 307 -240
rect 307 -241 308 -240
rect 308 -241 309 -240
rect 309 -241 310 -240
rect 310 -241 311 -240
rect 311 -241 312 -240
rect 312 -241 313 -240
rect 313 -241 314 -240
rect 314 -241 315 -240
rect 315 -241 316 -240
rect 316 -241 317 -240
rect 317 -241 318 -240
rect 318 -241 319 -240
rect 319 -241 320 -240
rect 320 -241 321 -240
rect 321 -241 322 -240
rect 322 -241 323 -240
rect 323 -241 324 -240
rect 324 -241 325 -240
rect 325 -241 326 -240
rect 326 -241 327 -240
rect 327 -241 328 -240
rect 328 -241 329 -240
rect 329 -241 330 -240
rect 330 -241 331 -240
rect 331 -241 332 -240
rect 332 -241 333 -240
rect 333 -241 334 -240
rect 334 -241 335 -240
rect 335 -241 336 -240
rect 336 -241 337 -240
rect 337 -241 338 -240
rect 338 -241 339 -240
rect 339 -241 340 -240
rect 340 -241 341 -240
rect 341 -241 342 -240
rect 342 -241 343 -240
rect 343 -241 344 -240
rect 344 -241 345 -240
rect 345 -241 346 -240
rect 346 -241 347 -240
rect 347 -241 348 -240
rect 348 -241 349 -240
rect 349 -241 350 -240
rect 350 -241 351 -240
rect 351 -241 352 -240
rect 352 -241 353 -240
rect 353 -241 354 -240
rect 354 -241 355 -240
rect 355 -241 356 -240
rect 356 -241 357 -240
rect 357 -241 358 -240
rect 358 -241 359 -240
rect 359 -241 360 -240
rect 360 -241 361 -240
rect 361 -241 362 -240
rect 362 -241 363 -240
rect 363 -241 364 -240
rect 364 -241 365 -240
rect 365 -241 366 -240
rect 366 -241 367 -240
rect 367 -241 368 -240
rect 368 -241 369 -240
rect 369 -241 370 -240
rect 370 -241 371 -240
rect 371 -241 372 -240
rect 372 -241 373 -240
rect 373 -241 374 -240
rect 374 -241 375 -240
rect 375 -241 376 -240
rect 376 -241 377 -240
rect 377 -241 378 -240
rect 378 -241 379 -240
rect 379 -241 380 -240
rect 380 -241 381 -240
rect 381 -241 382 -240
rect 382 -241 383 -240
rect 383 -241 384 -240
rect 384 -241 385 -240
rect 385 -241 386 -240
rect 386 -241 387 -240
rect 387 -241 388 -240
rect 388 -241 389 -240
rect 389 -241 390 -240
rect 390 -241 391 -240
rect 391 -241 392 -240
rect 392 -241 393 -240
rect 393 -241 394 -240
rect 394 -241 395 -240
rect 395 -241 396 -240
rect 396 -241 397 -240
rect 397 -241 398 -240
rect 398 -241 399 -240
rect 399 -241 400 -240
rect 400 -241 401 -240
rect 401 -241 402 -240
rect 402 -241 403 -240
rect 403 -241 404 -240
rect 404 -241 405 -240
rect 405 -241 406 -240
rect 406 -241 407 -240
rect 407 -241 408 -240
rect 408 -241 409 -240
rect 409 -241 410 -240
rect 410 -241 411 -240
rect 411 -241 412 -240
rect 412 -241 413 -240
rect 413 -241 414 -240
rect 414 -241 415 -240
rect 415 -241 416 -240
rect 416 -241 417 -240
rect 417 -241 418 -240
rect 418 -241 419 -240
rect 419 -241 420 -240
rect 420 -241 421 -240
rect 421 -241 422 -240
rect 422 -241 423 -240
rect 423 -241 424 -240
rect 424 -241 425 -240
rect 425 -241 426 -240
rect 426 -241 427 -240
rect 427 -241 428 -240
rect 428 -241 429 -240
rect 429 -241 430 -240
rect 430 -241 431 -240
rect 431 -241 432 -240
rect 432 -241 433 -240
rect 433 -241 434 -240
rect 434 -241 435 -240
rect 435 -241 436 -240
rect 436 -241 437 -240
rect 437 -241 438 -240
rect 438 -241 439 -240
rect 439 -241 440 -240
rect 440 -241 441 -240
rect 441 -241 442 -240
rect 442 -241 443 -240
rect 443 -241 444 -240
rect 444 -241 445 -240
rect 445 -241 446 -240
rect 446 -241 447 -240
rect 447 -241 448 -240
rect 448 -241 449 -240
rect 449 -241 450 -240
rect 450 -241 451 -240
rect 451 -241 452 -240
rect 452 -241 453 -240
rect 453 -241 454 -240
rect 454 -241 455 -240
rect 455 -241 456 -240
rect 456 -241 457 -240
rect 457 -241 458 -240
rect 458 -241 459 -240
rect 459 -241 460 -240
rect 460 -241 461 -240
rect 461 -241 462 -240
rect 462 -241 463 -240
rect 463 -241 464 -240
rect 464 -241 465 -240
rect 465 -241 466 -240
rect 466 -241 467 -240
rect 467 -241 468 -240
rect 468 -241 469 -240
rect 469 -241 470 -240
rect 470 -241 471 -240
rect 471 -241 472 -240
rect 472 -241 473 -240
rect 473 -241 474 -240
rect 474 -241 475 -240
rect 475 -241 476 -240
rect 476 -241 477 -240
rect 477 -241 478 -240
rect 478 -241 479 -240
rect 479 -241 480 -240
rect 2 -242 3 -241
rect 3 -242 4 -241
rect 4 -242 5 -241
rect 5 -242 6 -241
rect 6 -242 7 -241
rect 7 -242 8 -241
rect 8 -242 9 -241
rect 9 -242 10 -241
rect 10 -242 11 -241
rect 11 -242 12 -241
rect 12 -242 13 -241
rect 13 -242 14 -241
rect 14 -242 15 -241
rect 15 -242 16 -241
rect 16 -242 17 -241
rect 17 -242 18 -241
rect 18 -242 19 -241
rect 19 -242 20 -241
rect 20 -242 21 -241
rect 21 -242 22 -241
rect 22 -242 23 -241
rect 23 -242 24 -241
rect 24 -242 25 -241
rect 25 -242 26 -241
rect 26 -242 27 -241
rect 27 -242 28 -241
rect 28 -242 29 -241
rect 29 -242 30 -241
rect 30 -242 31 -241
rect 31 -242 32 -241
rect 32 -242 33 -241
rect 33 -242 34 -241
rect 34 -242 35 -241
rect 35 -242 36 -241
rect 36 -242 37 -241
rect 37 -242 38 -241
rect 38 -242 39 -241
rect 39 -242 40 -241
rect 40 -242 41 -241
rect 41 -242 42 -241
rect 42 -242 43 -241
rect 43 -242 44 -241
rect 44 -242 45 -241
rect 45 -242 46 -241
rect 46 -242 47 -241
rect 47 -242 48 -241
rect 48 -242 49 -241
rect 49 -242 50 -241
rect 50 -242 51 -241
rect 51 -242 52 -241
rect 52 -242 53 -241
rect 53 -242 54 -241
rect 54 -242 55 -241
rect 55 -242 56 -241
rect 56 -242 57 -241
rect 57 -242 58 -241
rect 58 -242 59 -241
rect 59 -242 60 -241
rect 60 -242 61 -241
rect 61 -242 62 -241
rect 62 -242 63 -241
rect 63 -242 64 -241
rect 64 -242 65 -241
rect 65 -242 66 -241
rect 66 -242 67 -241
rect 67 -242 68 -241
rect 68 -242 69 -241
rect 69 -242 70 -241
rect 70 -242 71 -241
rect 71 -242 72 -241
rect 72 -242 73 -241
rect 73 -242 74 -241
rect 74 -242 75 -241
rect 75 -242 76 -241
rect 76 -242 77 -241
rect 77 -242 78 -241
rect 78 -242 79 -241
rect 79 -242 80 -241
rect 80 -242 81 -241
rect 81 -242 82 -241
rect 82 -242 83 -241
rect 83 -242 84 -241
rect 84 -242 85 -241
rect 85 -242 86 -241
rect 86 -242 87 -241
rect 87 -242 88 -241
rect 88 -242 89 -241
rect 89 -242 90 -241
rect 90 -242 91 -241
rect 91 -242 92 -241
rect 92 -242 93 -241
rect 93 -242 94 -241
rect 94 -242 95 -241
rect 95 -242 96 -241
rect 96 -242 97 -241
rect 97 -242 98 -241
rect 98 -242 99 -241
rect 99 -242 100 -241
rect 100 -242 101 -241
rect 101 -242 102 -241
rect 102 -242 103 -241
rect 103 -242 104 -241
rect 104 -242 105 -241
rect 105 -242 106 -241
rect 106 -242 107 -241
rect 107 -242 108 -241
rect 108 -242 109 -241
rect 109 -242 110 -241
rect 110 -242 111 -241
rect 111 -242 112 -241
rect 112 -242 113 -241
rect 113 -242 114 -241
rect 114 -242 115 -241
rect 115 -242 116 -241
rect 116 -242 117 -241
rect 117 -242 118 -241
rect 118 -242 119 -241
rect 119 -242 120 -241
rect 120 -242 121 -241
rect 121 -242 122 -241
rect 122 -242 123 -241
rect 123 -242 124 -241
rect 124 -242 125 -241
rect 125 -242 126 -241
rect 126 -242 127 -241
rect 127 -242 128 -241
rect 128 -242 129 -241
rect 129 -242 130 -241
rect 130 -242 131 -241
rect 131 -242 132 -241
rect 132 -242 133 -241
rect 133 -242 134 -241
rect 134 -242 135 -241
rect 135 -242 136 -241
rect 136 -242 137 -241
rect 137 -242 138 -241
rect 138 -242 139 -241
rect 139 -242 140 -241
rect 140 -242 141 -241
rect 141 -242 142 -241
rect 142 -242 143 -241
rect 143 -242 144 -241
rect 144 -242 145 -241
rect 145 -242 146 -241
rect 146 -242 147 -241
rect 147 -242 148 -241
rect 148 -242 149 -241
rect 149 -242 150 -241
rect 150 -242 151 -241
rect 151 -242 152 -241
rect 152 -242 153 -241
rect 153 -242 154 -241
rect 154 -242 155 -241
rect 155 -242 156 -241
rect 156 -242 157 -241
rect 157 -242 158 -241
rect 158 -242 159 -241
rect 159 -242 160 -241
rect 160 -242 161 -241
rect 161 -242 162 -241
rect 162 -242 163 -241
rect 163 -242 164 -241
rect 164 -242 165 -241
rect 165 -242 166 -241
rect 166 -242 167 -241
rect 167 -242 168 -241
rect 168 -242 169 -241
rect 169 -242 170 -241
rect 170 -242 171 -241
rect 171 -242 172 -241
rect 172 -242 173 -241
rect 173 -242 174 -241
rect 174 -242 175 -241
rect 175 -242 176 -241
rect 176 -242 177 -241
rect 177 -242 178 -241
rect 178 -242 179 -241
rect 179 -242 180 -241
rect 180 -242 181 -241
rect 181 -242 182 -241
rect 182 -242 183 -241
rect 183 -242 184 -241
rect 184 -242 185 -241
rect 185 -242 186 -241
rect 186 -242 187 -241
rect 187 -242 188 -241
rect 188 -242 189 -241
rect 189 -242 190 -241
rect 190 -242 191 -241
rect 191 -242 192 -241
rect 192 -242 193 -241
rect 193 -242 194 -241
rect 194 -242 195 -241
rect 195 -242 196 -241
rect 196 -242 197 -241
rect 197 -242 198 -241
rect 198 -242 199 -241
rect 199 -242 200 -241
rect 200 -242 201 -241
rect 201 -242 202 -241
rect 202 -242 203 -241
rect 203 -242 204 -241
rect 204 -242 205 -241
rect 205 -242 206 -241
rect 206 -242 207 -241
rect 207 -242 208 -241
rect 208 -242 209 -241
rect 209 -242 210 -241
rect 210 -242 211 -241
rect 211 -242 212 -241
rect 212 -242 213 -241
rect 213 -242 214 -241
rect 214 -242 215 -241
rect 215 -242 216 -241
rect 216 -242 217 -241
rect 217 -242 218 -241
rect 218 -242 219 -241
rect 219 -242 220 -241
rect 220 -242 221 -241
rect 221 -242 222 -241
rect 222 -242 223 -241
rect 223 -242 224 -241
rect 224 -242 225 -241
rect 225 -242 226 -241
rect 226 -242 227 -241
rect 227 -242 228 -241
rect 228 -242 229 -241
rect 229 -242 230 -241
rect 230 -242 231 -241
rect 231 -242 232 -241
rect 232 -242 233 -241
rect 233 -242 234 -241
rect 234 -242 235 -241
rect 235 -242 236 -241
rect 236 -242 237 -241
rect 237 -242 238 -241
rect 238 -242 239 -241
rect 239 -242 240 -241
rect 240 -242 241 -241
rect 241 -242 242 -241
rect 242 -242 243 -241
rect 243 -242 244 -241
rect 244 -242 245 -241
rect 245 -242 246 -241
rect 246 -242 247 -241
rect 247 -242 248 -241
rect 248 -242 249 -241
rect 249 -242 250 -241
rect 250 -242 251 -241
rect 251 -242 252 -241
rect 252 -242 253 -241
rect 253 -242 254 -241
rect 254 -242 255 -241
rect 255 -242 256 -241
rect 256 -242 257 -241
rect 257 -242 258 -241
rect 258 -242 259 -241
rect 259 -242 260 -241
rect 260 -242 261 -241
rect 261 -242 262 -241
rect 262 -242 263 -241
rect 263 -242 264 -241
rect 264 -242 265 -241
rect 265 -242 266 -241
rect 266 -242 267 -241
rect 267 -242 268 -241
rect 268 -242 269 -241
rect 269 -242 270 -241
rect 270 -242 271 -241
rect 271 -242 272 -241
rect 272 -242 273 -241
rect 273 -242 274 -241
rect 274 -242 275 -241
rect 275 -242 276 -241
rect 276 -242 277 -241
rect 277 -242 278 -241
rect 278 -242 279 -241
rect 279 -242 280 -241
rect 280 -242 281 -241
rect 281 -242 282 -241
rect 282 -242 283 -241
rect 283 -242 284 -241
rect 284 -242 285 -241
rect 285 -242 286 -241
rect 286 -242 287 -241
rect 287 -242 288 -241
rect 288 -242 289 -241
rect 289 -242 290 -241
rect 290 -242 291 -241
rect 291 -242 292 -241
rect 292 -242 293 -241
rect 293 -242 294 -241
rect 294 -242 295 -241
rect 295 -242 296 -241
rect 296 -242 297 -241
rect 297 -242 298 -241
rect 298 -242 299 -241
rect 299 -242 300 -241
rect 300 -242 301 -241
rect 301 -242 302 -241
rect 302 -242 303 -241
rect 303 -242 304 -241
rect 304 -242 305 -241
rect 305 -242 306 -241
rect 306 -242 307 -241
rect 307 -242 308 -241
rect 308 -242 309 -241
rect 309 -242 310 -241
rect 310 -242 311 -241
rect 311 -242 312 -241
rect 312 -242 313 -241
rect 313 -242 314 -241
rect 314 -242 315 -241
rect 315 -242 316 -241
rect 316 -242 317 -241
rect 317 -242 318 -241
rect 318 -242 319 -241
rect 319 -242 320 -241
rect 320 -242 321 -241
rect 321 -242 322 -241
rect 322 -242 323 -241
rect 323 -242 324 -241
rect 324 -242 325 -241
rect 325 -242 326 -241
rect 326 -242 327 -241
rect 327 -242 328 -241
rect 328 -242 329 -241
rect 329 -242 330 -241
rect 330 -242 331 -241
rect 331 -242 332 -241
rect 332 -242 333 -241
rect 333 -242 334 -241
rect 334 -242 335 -241
rect 335 -242 336 -241
rect 336 -242 337 -241
rect 337 -242 338 -241
rect 338 -242 339 -241
rect 339 -242 340 -241
rect 340 -242 341 -241
rect 341 -242 342 -241
rect 342 -242 343 -241
rect 343 -242 344 -241
rect 344 -242 345 -241
rect 345 -242 346 -241
rect 346 -242 347 -241
rect 347 -242 348 -241
rect 348 -242 349 -241
rect 349 -242 350 -241
rect 350 -242 351 -241
rect 351 -242 352 -241
rect 352 -242 353 -241
rect 353 -242 354 -241
rect 354 -242 355 -241
rect 355 -242 356 -241
rect 356 -242 357 -241
rect 357 -242 358 -241
rect 358 -242 359 -241
rect 359 -242 360 -241
rect 360 -242 361 -241
rect 361 -242 362 -241
rect 362 -242 363 -241
rect 363 -242 364 -241
rect 364 -242 365 -241
rect 365 -242 366 -241
rect 366 -242 367 -241
rect 367 -242 368 -241
rect 368 -242 369 -241
rect 369 -242 370 -241
rect 370 -242 371 -241
rect 371 -242 372 -241
rect 372 -242 373 -241
rect 373 -242 374 -241
rect 374 -242 375 -241
rect 375 -242 376 -241
rect 376 -242 377 -241
rect 377 -242 378 -241
rect 378 -242 379 -241
rect 379 -242 380 -241
rect 380 -242 381 -241
rect 381 -242 382 -241
rect 382 -242 383 -241
rect 383 -242 384 -241
rect 384 -242 385 -241
rect 385 -242 386 -241
rect 386 -242 387 -241
rect 387 -242 388 -241
rect 388 -242 389 -241
rect 389 -242 390 -241
rect 390 -242 391 -241
rect 391 -242 392 -241
rect 392 -242 393 -241
rect 393 -242 394 -241
rect 394 -242 395 -241
rect 395 -242 396 -241
rect 396 -242 397 -241
rect 397 -242 398 -241
rect 398 -242 399 -241
rect 399 -242 400 -241
rect 400 -242 401 -241
rect 401 -242 402 -241
rect 402 -242 403 -241
rect 403 -242 404 -241
rect 404 -242 405 -241
rect 405 -242 406 -241
rect 406 -242 407 -241
rect 407 -242 408 -241
rect 408 -242 409 -241
rect 409 -242 410 -241
rect 410 -242 411 -241
rect 411 -242 412 -241
rect 412 -242 413 -241
rect 413 -242 414 -241
rect 414 -242 415 -241
rect 415 -242 416 -241
rect 416 -242 417 -241
rect 417 -242 418 -241
rect 418 -242 419 -241
rect 419 -242 420 -241
rect 420 -242 421 -241
rect 421 -242 422 -241
rect 422 -242 423 -241
rect 423 -242 424 -241
rect 424 -242 425 -241
rect 425 -242 426 -241
rect 426 -242 427 -241
rect 427 -242 428 -241
rect 428 -242 429 -241
rect 429 -242 430 -241
rect 430 -242 431 -241
rect 431 -242 432 -241
rect 432 -242 433 -241
rect 433 -242 434 -241
rect 434 -242 435 -241
rect 435 -242 436 -241
rect 436 -242 437 -241
rect 437 -242 438 -241
rect 438 -242 439 -241
rect 439 -242 440 -241
rect 440 -242 441 -241
rect 441 -242 442 -241
rect 442 -242 443 -241
rect 443 -242 444 -241
rect 444 -242 445 -241
rect 445 -242 446 -241
rect 446 -242 447 -241
rect 447 -242 448 -241
rect 448 -242 449 -241
rect 449 -242 450 -241
rect 450 -242 451 -241
rect 451 -242 452 -241
rect 452 -242 453 -241
rect 453 -242 454 -241
rect 454 -242 455 -241
rect 455 -242 456 -241
rect 456 -242 457 -241
rect 457 -242 458 -241
rect 458 -242 459 -241
rect 459 -242 460 -241
rect 460 -242 461 -241
rect 461 -242 462 -241
rect 462 -242 463 -241
rect 463 -242 464 -241
rect 464 -242 465 -241
rect 465 -242 466 -241
rect 466 -242 467 -241
rect 467 -242 468 -241
rect 468 -242 469 -241
rect 469 -242 470 -241
rect 470 -242 471 -241
rect 471 -242 472 -241
rect 472 -242 473 -241
rect 473 -242 474 -241
rect 474 -242 475 -241
rect 475 -242 476 -241
rect 476 -242 477 -241
rect 477 -242 478 -241
rect 478 -242 479 -241
rect 479 -242 480 -241
rect 2 -243 3 -242
rect 3 -243 4 -242
rect 4 -243 5 -242
rect 5 -243 6 -242
rect 6 -243 7 -242
rect 7 -243 8 -242
rect 8 -243 9 -242
rect 9 -243 10 -242
rect 10 -243 11 -242
rect 11 -243 12 -242
rect 12 -243 13 -242
rect 13 -243 14 -242
rect 14 -243 15 -242
rect 15 -243 16 -242
rect 16 -243 17 -242
rect 17 -243 18 -242
rect 18 -243 19 -242
rect 19 -243 20 -242
rect 20 -243 21 -242
rect 21 -243 22 -242
rect 22 -243 23 -242
rect 23 -243 24 -242
rect 24 -243 25 -242
rect 25 -243 26 -242
rect 26 -243 27 -242
rect 27 -243 28 -242
rect 28 -243 29 -242
rect 29 -243 30 -242
rect 30 -243 31 -242
rect 31 -243 32 -242
rect 32 -243 33 -242
rect 33 -243 34 -242
rect 34 -243 35 -242
rect 35 -243 36 -242
rect 36 -243 37 -242
rect 37 -243 38 -242
rect 38 -243 39 -242
rect 39 -243 40 -242
rect 40 -243 41 -242
rect 41 -243 42 -242
rect 42 -243 43 -242
rect 43 -243 44 -242
rect 44 -243 45 -242
rect 45 -243 46 -242
rect 46 -243 47 -242
rect 47 -243 48 -242
rect 48 -243 49 -242
rect 49 -243 50 -242
rect 50 -243 51 -242
rect 51 -243 52 -242
rect 52 -243 53 -242
rect 53 -243 54 -242
rect 54 -243 55 -242
rect 55 -243 56 -242
rect 56 -243 57 -242
rect 57 -243 58 -242
rect 58 -243 59 -242
rect 59 -243 60 -242
rect 60 -243 61 -242
rect 61 -243 62 -242
rect 62 -243 63 -242
rect 63 -243 64 -242
rect 64 -243 65 -242
rect 65 -243 66 -242
rect 66 -243 67 -242
rect 67 -243 68 -242
rect 68 -243 69 -242
rect 69 -243 70 -242
rect 70 -243 71 -242
rect 71 -243 72 -242
rect 72 -243 73 -242
rect 73 -243 74 -242
rect 74 -243 75 -242
rect 75 -243 76 -242
rect 76 -243 77 -242
rect 77 -243 78 -242
rect 78 -243 79 -242
rect 79 -243 80 -242
rect 80 -243 81 -242
rect 81 -243 82 -242
rect 82 -243 83 -242
rect 83 -243 84 -242
rect 84 -243 85 -242
rect 85 -243 86 -242
rect 86 -243 87 -242
rect 87 -243 88 -242
rect 88 -243 89 -242
rect 89 -243 90 -242
rect 90 -243 91 -242
rect 91 -243 92 -242
rect 92 -243 93 -242
rect 93 -243 94 -242
rect 94 -243 95 -242
rect 95 -243 96 -242
rect 96 -243 97 -242
rect 97 -243 98 -242
rect 98 -243 99 -242
rect 99 -243 100 -242
rect 100 -243 101 -242
rect 101 -243 102 -242
rect 102 -243 103 -242
rect 103 -243 104 -242
rect 104 -243 105 -242
rect 105 -243 106 -242
rect 106 -243 107 -242
rect 107 -243 108 -242
rect 108 -243 109 -242
rect 109 -243 110 -242
rect 110 -243 111 -242
rect 111 -243 112 -242
rect 112 -243 113 -242
rect 113 -243 114 -242
rect 114 -243 115 -242
rect 115 -243 116 -242
rect 116 -243 117 -242
rect 117 -243 118 -242
rect 118 -243 119 -242
rect 119 -243 120 -242
rect 120 -243 121 -242
rect 121 -243 122 -242
rect 122 -243 123 -242
rect 123 -243 124 -242
rect 124 -243 125 -242
rect 125 -243 126 -242
rect 126 -243 127 -242
rect 127 -243 128 -242
rect 128 -243 129 -242
rect 129 -243 130 -242
rect 130 -243 131 -242
rect 131 -243 132 -242
rect 132 -243 133 -242
rect 133 -243 134 -242
rect 134 -243 135 -242
rect 135 -243 136 -242
rect 136 -243 137 -242
rect 137 -243 138 -242
rect 138 -243 139 -242
rect 139 -243 140 -242
rect 140 -243 141 -242
rect 141 -243 142 -242
rect 142 -243 143 -242
rect 143 -243 144 -242
rect 144 -243 145 -242
rect 145 -243 146 -242
rect 146 -243 147 -242
rect 147 -243 148 -242
rect 148 -243 149 -242
rect 149 -243 150 -242
rect 150 -243 151 -242
rect 151 -243 152 -242
rect 152 -243 153 -242
rect 153 -243 154 -242
rect 154 -243 155 -242
rect 155 -243 156 -242
rect 156 -243 157 -242
rect 157 -243 158 -242
rect 158 -243 159 -242
rect 159 -243 160 -242
rect 160 -243 161 -242
rect 161 -243 162 -242
rect 162 -243 163 -242
rect 163 -243 164 -242
rect 164 -243 165 -242
rect 165 -243 166 -242
rect 166 -243 167 -242
rect 167 -243 168 -242
rect 168 -243 169 -242
rect 169 -243 170 -242
rect 170 -243 171 -242
rect 171 -243 172 -242
rect 172 -243 173 -242
rect 173 -243 174 -242
rect 174 -243 175 -242
rect 175 -243 176 -242
rect 176 -243 177 -242
rect 177 -243 178 -242
rect 178 -243 179 -242
rect 179 -243 180 -242
rect 180 -243 181 -242
rect 181 -243 182 -242
rect 182 -243 183 -242
rect 183 -243 184 -242
rect 184 -243 185 -242
rect 185 -243 186 -242
rect 186 -243 187 -242
rect 187 -243 188 -242
rect 188 -243 189 -242
rect 189 -243 190 -242
rect 190 -243 191 -242
rect 191 -243 192 -242
rect 192 -243 193 -242
rect 193 -243 194 -242
rect 194 -243 195 -242
rect 195 -243 196 -242
rect 196 -243 197 -242
rect 197 -243 198 -242
rect 198 -243 199 -242
rect 199 -243 200 -242
rect 200 -243 201 -242
rect 201 -243 202 -242
rect 202 -243 203 -242
rect 203 -243 204 -242
rect 204 -243 205 -242
rect 205 -243 206 -242
rect 206 -243 207 -242
rect 207 -243 208 -242
rect 208 -243 209 -242
rect 209 -243 210 -242
rect 210 -243 211 -242
rect 211 -243 212 -242
rect 212 -243 213 -242
rect 213 -243 214 -242
rect 214 -243 215 -242
rect 215 -243 216 -242
rect 216 -243 217 -242
rect 217 -243 218 -242
rect 218 -243 219 -242
rect 219 -243 220 -242
rect 220 -243 221 -242
rect 221 -243 222 -242
rect 222 -243 223 -242
rect 223 -243 224 -242
rect 224 -243 225 -242
rect 225 -243 226 -242
rect 226 -243 227 -242
rect 227 -243 228 -242
rect 228 -243 229 -242
rect 229 -243 230 -242
rect 230 -243 231 -242
rect 231 -243 232 -242
rect 232 -243 233 -242
rect 233 -243 234 -242
rect 234 -243 235 -242
rect 235 -243 236 -242
rect 236 -243 237 -242
rect 237 -243 238 -242
rect 238 -243 239 -242
rect 239 -243 240 -242
rect 240 -243 241 -242
rect 241 -243 242 -242
rect 242 -243 243 -242
rect 243 -243 244 -242
rect 244 -243 245 -242
rect 245 -243 246 -242
rect 246 -243 247 -242
rect 247 -243 248 -242
rect 248 -243 249 -242
rect 249 -243 250 -242
rect 250 -243 251 -242
rect 251 -243 252 -242
rect 252 -243 253 -242
rect 253 -243 254 -242
rect 254 -243 255 -242
rect 255 -243 256 -242
rect 256 -243 257 -242
rect 257 -243 258 -242
rect 258 -243 259 -242
rect 259 -243 260 -242
rect 260 -243 261 -242
rect 261 -243 262 -242
rect 262 -243 263 -242
rect 263 -243 264 -242
rect 264 -243 265 -242
rect 265 -243 266 -242
rect 266 -243 267 -242
rect 267 -243 268 -242
rect 268 -243 269 -242
rect 269 -243 270 -242
rect 270 -243 271 -242
rect 271 -243 272 -242
rect 272 -243 273 -242
rect 273 -243 274 -242
rect 274 -243 275 -242
rect 275 -243 276 -242
rect 276 -243 277 -242
rect 277 -243 278 -242
rect 278 -243 279 -242
rect 279 -243 280 -242
rect 280 -243 281 -242
rect 281 -243 282 -242
rect 282 -243 283 -242
rect 283 -243 284 -242
rect 284 -243 285 -242
rect 285 -243 286 -242
rect 286 -243 287 -242
rect 287 -243 288 -242
rect 288 -243 289 -242
rect 289 -243 290 -242
rect 290 -243 291 -242
rect 291 -243 292 -242
rect 292 -243 293 -242
rect 293 -243 294 -242
rect 294 -243 295 -242
rect 295 -243 296 -242
rect 296 -243 297 -242
rect 297 -243 298 -242
rect 298 -243 299 -242
rect 299 -243 300 -242
rect 300 -243 301 -242
rect 301 -243 302 -242
rect 302 -243 303 -242
rect 303 -243 304 -242
rect 304 -243 305 -242
rect 305 -243 306 -242
rect 306 -243 307 -242
rect 307 -243 308 -242
rect 308 -243 309 -242
rect 309 -243 310 -242
rect 310 -243 311 -242
rect 311 -243 312 -242
rect 312 -243 313 -242
rect 313 -243 314 -242
rect 314 -243 315 -242
rect 315 -243 316 -242
rect 316 -243 317 -242
rect 317 -243 318 -242
rect 318 -243 319 -242
rect 319 -243 320 -242
rect 320 -243 321 -242
rect 321 -243 322 -242
rect 322 -243 323 -242
rect 323 -243 324 -242
rect 324 -243 325 -242
rect 325 -243 326 -242
rect 326 -243 327 -242
rect 327 -243 328 -242
rect 328 -243 329 -242
rect 329 -243 330 -242
rect 330 -243 331 -242
rect 331 -243 332 -242
rect 332 -243 333 -242
rect 333 -243 334 -242
rect 334 -243 335 -242
rect 335 -243 336 -242
rect 336 -243 337 -242
rect 337 -243 338 -242
rect 338 -243 339 -242
rect 339 -243 340 -242
rect 340 -243 341 -242
rect 341 -243 342 -242
rect 342 -243 343 -242
rect 343 -243 344 -242
rect 344 -243 345 -242
rect 345 -243 346 -242
rect 346 -243 347 -242
rect 347 -243 348 -242
rect 348 -243 349 -242
rect 349 -243 350 -242
rect 350 -243 351 -242
rect 351 -243 352 -242
rect 352 -243 353 -242
rect 353 -243 354 -242
rect 354 -243 355 -242
rect 355 -243 356 -242
rect 356 -243 357 -242
rect 357 -243 358 -242
rect 358 -243 359 -242
rect 359 -243 360 -242
rect 360 -243 361 -242
rect 361 -243 362 -242
rect 362 -243 363 -242
rect 363 -243 364 -242
rect 364 -243 365 -242
rect 365 -243 366 -242
rect 366 -243 367 -242
rect 367 -243 368 -242
rect 368 -243 369 -242
rect 369 -243 370 -242
rect 370 -243 371 -242
rect 371 -243 372 -242
rect 372 -243 373 -242
rect 373 -243 374 -242
rect 374 -243 375 -242
rect 375 -243 376 -242
rect 376 -243 377 -242
rect 377 -243 378 -242
rect 378 -243 379 -242
rect 379 -243 380 -242
rect 380 -243 381 -242
rect 381 -243 382 -242
rect 382 -243 383 -242
rect 383 -243 384 -242
rect 384 -243 385 -242
rect 385 -243 386 -242
rect 386 -243 387 -242
rect 387 -243 388 -242
rect 388 -243 389 -242
rect 389 -243 390 -242
rect 390 -243 391 -242
rect 391 -243 392 -242
rect 392 -243 393 -242
rect 393 -243 394 -242
rect 394 -243 395 -242
rect 395 -243 396 -242
rect 396 -243 397 -242
rect 397 -243 398 -242
rect 398 -243 399 -242
rect 399 -243 400 -242
rect 400 -243 401 -242
rect 401 -243 402 -242
rect 402 -243 403 -242
rect 403 -243 404 -242
rect 404 -243 405 -242
rect 405 -243 406 -242
rect 406 -243 407 -242
rect 407 -243 408 -242
rect 408 -243 409 -242
rect 409 -243 410 -242
rect 410 -243 411 -242
rect 411 -243 412 -242
rect 412 -243 413 -242
rect 413 -243 414 -242
rect 414 -243 415 -242
rect 415 -243 416 -242
rect 416 -243 417 -242
rect 417 -243 418 -242
rect 418 -243 419 -242
rect 419 -243 420 -242
rect 420 -243 421 -242
rect 421 -243 422 -242
rect 422 -243 423 -242
rect 423 -243 424 -242
rect 424 -243 425 -242
rect 425 -243 426 -242
rect 426 -243 427 -242
rect 427 -243 428 -242
rect 428 -243 429 -242
rect 429 -243 430 -242
rect 430 -243 431 -242
rect 431 -243 432 -242
rect 432 -243 433 -242
rect 433 -243 434 -242
rect 434 -243 435 -242
rect 435 -243 436 -242
rect 436 -243 437 -242
rect 437 -243 438 -242
rect 438 -243 439 -242
rect 439 -243 440 -242
rect 440 -243 441 -242
rect 441 -243 442 -242
rect 442 -243 443 -242
rect 443 -243 444 -242
rect 444 -243 445 -242
rect 445 -243 446 -242
rect 446 -243 447 -242
rect 447 -243 448 -242
rect 448 -243 449 -242
rect 449 -243 450 -242
rect 450 -243 451 -242
rect 451 -243 452 -242
rect 452 -243 453 -242
rect 453 -243 454 -242
rect 454 -243 455 -242
rect 455 -243 456 -242
rect 456 -243 457 -242
rect 457 -243 458 -242
rect 458 -243 459 -242
rect 459 -243 460 -242
rect 460 -243 461 -242
rect 461 -243 462 -242
rect 462 -243 463 -242
rect 463 -243 464 -242
rect 464 -243 465 -242
rect 465 -243 466 -242
rect 466 -243 467 -242
rect 467 -243 468 -242
rect 468 -243 469 -242
rect 469 -243 470 -242
rect 470 -243 471 -242
rect 471 -243 472 -242
rect 472 -243 473 -242
rect 473 -243 474 -242
rect 474 -243 475 -242
rect 475 -243 476 -242
rect 476 -243 477 -242
rect 477 -243 478 -242
rect 478 -243 479 -242
rect 479 -243 480 -242
rect 2 -244 3 -243
rect 3 -244 4 -243
rect 4 -244 5 -243
rect 5 -244 6 -243
rect 6 -244 7 -243
rect 7 -244 8 -243
rect 8 -244 9 -243
rect 9 -244 10 -243
rect 10 -244 11 -243
rect 11 -244 12 -243
rect 12 -244 13 -243
rect 13 -244 14 -243
rect 14 -244 15 -243
rect 15 -244 16 -243
rect 16 -244 17 -243
rect 17 -244 18 -243
rect 18 -244 19 -243
rect 19 -244 20 -243
rect 20 -244 21 -243
rect 21 -244 22 -243
rect 22 -244 23 -243
rect 23 -244 24 -243
rect 24 -244 25 -243
rect 25 -244 26 -243
rect 26 -244 27 -243
rect 27 -244 28 -243
rect 28 -244 29 -243
rect 29 -244 30 -243
rect 30 -244 31 -243
rect 31 -244 32 -243
rect 32 -244 33 -243
rect 33 -244 34 -243
rect 34 -244 35 -243
rect 35 -244 36 -243
rect 36 -244 37 -243
rect 37 -244 38 -243
rect 38 -244 39 -243
rect 39 -244 40 -243
rect 40 -244 41 -243
rect 41 -244 42 -243
rect 42 -244 43 -243
rect 43 -244 44 -243
rect 44 -244 45 -243
rect 45 -244 46 -243
rect 46 -244 47 -243
rect 47 -244 48 -243
rect 48 -244 49 -243
rect 49 -244 50 -243
rect 50 -244 51 -243
rect 51 -244 52 -243
rect 52 -244 53 -243
rect 53 -244 54 -243
rect 54 -244 55 -243
rect 55 -244 56 -243
rect 56 -244 57 -243
rect 57 -244 58 -243
rect 58 -244 59 -243
rect 59 -244 60 -243
rect 60 -244 61 -243
rect 61 -244 62 -243
rect 62 -244 63 -243
rect 63 -244 64 -243
rect 64 -244 65 -243
rect 65 -244 66 -243
rect 66 -244 67 -243
rect 67 -244 68 -243
rect 68 -244 69 -243
rect 69 -244 70 -243
rect 70 -244 71 -243
rect 71 -244 72 -243
rect 72 -244 73 -243
rect 73 -244 74 -243
rect 74 -244 75 -243
rect 75 -244 76 -243
rect 76 -244 77 -243
rect 77 -244 78 -243
rect 78 -244 79 -243
rect 79 -244 80 -243
rect 80 -244 81 -243
rect 81 -244 82 -243
rect 82 -244 83 -243
rect 83 -244 84 -243
rect 84 -244 85 -243
rect 85 -244 86 -243
rect 86 -244 87 -243
rect 87 -244 88 -243
rect 88 -244 89 -243
rect 89 -244 90 -243
rect 90 -244 91 -243
rect 91 -244 92 -243
rect 92 -244 93 -243
rect 93 -244 94 -243
rect 94 -244 95 -243
rect 95 -244 96 -243
rect 96 -244 97 -243
rect 97 -244 98 -243
rect 98 -244 99 -243
rect 99 -244 100 -243
rect 100 -244 101 -243
rect 101 -244 102 -243
rect 102 -244 103 -243
rect 103 -244 104 -243
rect 104 -244 105 -243
rect 105 -244 106 -243
rect 106 -244 107 -243
rect 107 -244 108 -243
rect 108 -244 109 -243
rect 109 -244 110 -243
rect 110 -244 111 -243
rect 111 -244 112 -243
rect 112 -244 113 -243
rect 113 -244 114 -243
rect 114 -244 115 -243
rect 115 -244 116 -243
rect 116 -244 117 -243
rect 117 -244 118 -243
rect 118 -244 119 -243
rect 119 -244 120 -243
rect 120 -244 121 -243
rect 121 -244 122 -243
rect 122 -244 123 -243
rect 123 -244 124 -243
rect 124 -244 125 -243
rect 125 -244 126 -243
rect 126 -244 127 -243
rect 127 -244 128 -243
rect 128 -244 129 -243
rect 129 -244 130 -243
rect 130 -244 131 -243
rect 131 -244 132 -243
rect 132 -244 133 -243
rect 133 -244 134 -243
rect 134 -244 135 -243
rect 135 -244 136 -243
rect 136 -244 137 -243
rect 137 -244 138 -243
rect 138 -244 139 -243
rect 139 -244 140 -243
rect 140 -244 141 -243
rect 141 -244 142 -243
rect 142 -244 143 -243
rect 143 -244 144 -243
rect 144 -244 145 -243
rect 145 -244 146 -243
rect 146 -244 147 -243
rect 147 -244 148 -243
rect 148 -244 149 -243
rect 149 -244 150 -243
rect 150 -244 151 -243
rect 151 -244 152 -243
rect 152 -244 153 -243
rect 153 -244 154 -243
rect 154 -244 155 -243
rect 155 -244 156 -243
rect 156 -244 157 -243
rect 157 -244 158 -243
rect 158 -244 159 -243
rect 159 -244 160 -243
rect 160 -244 161 -243
rect 161 -244 162 -243
rect 162 -244 163 -243
rect 163 -244 164 -243
rect 164 -244 165 -243
rect 165 -244 166 -243
rect 166 -244 167 -243
rect 167 -244 168 -243
rect 168 -244 169 -243
rect 169 -244 170 -243
rect 170 -244 171 -243
rect 171 -244 172 -243
rect 172 -244 173 -243
rect 173 -244 174 -243
rect 174 -244 175 -243
rect 175 -244 176 -243
rect 176 -244 177 -243
rect 177 -244 178 -243
rect 178 -244 179 -243
rect 179 -244 180 -243
rect 180 -244 181 -243
rect 181 -244 182 -243
rect 182 -244 183 -243
rect 183 -244 184 -243
rect 184 -244 185 -243
rect 185 -244 186 -243
rect 186 -244 187 -243
rect 187 -244 188 -243
rect 188 -244 189 -243
rect 189 -244 190 -243
rect 190 -244 191 -243
rect 191 -244 192 -243
rect 192 -244 193 -243
rect 193 -244 194 -243
rect 194 -244 195 -243
rect 195 -244 196 -243
rect 196 -244 197 -243
rect 197 -244 198 -243
rect 198 -244 199 -243
rect 199 -244 200 -243
rect 200 -244 201 -243
rect 201 -244 202 -243
rect 202 -244 203 -243
rect 203 -244 204 -243
rect 204 -244 205 -243
rect 205 -244 206 -243
rect 206 -244 207 -243
rect 207 -244 208 -243
rect 208 -244 209 -243
rect 209 -244 210 -243
rect 210 -244 211 -243
rect 211 -244 212 -243
rect 212 -244 213 -243
rect 213 -244 214 -243
rect 214 -244 215 -243
rect 215 -244 216 -243
rect 216 -244 217 -243
rect 217 -244 218 -243
rect 218 -244 219 -243
rect 219 -244 220 -243
rect 220 -244 221 -243
rect 221 -244 222 -243
rect 222 -244 223 -243
rect 223 -244 224 -243
rect 224 -244 225 -243
rect 225 -244 226 -243
rect 226 -244 227 -243
rect 227 -244 228 -243
rect 228 -244 229 -243
rect 229 -244 230 -243
rect 230 -244 231 -243
rect 231 -244 232 -243
rect 232 -244 233 -243
rect 233 -244 234 -243
rect 234 -244 235 -243
rect 235 -244 236 -243
rect 236 -244 237 -243
rect 237 -244 238 -243
rect 238 -244 239 -243
rect 239 -244 240 -243
rect 240 -244 241 -243
rect 241 -244 242 -243
rect 242 -244 243 -243
rect 243 -244 244 -243
rect 244 -244 245 -243
rect 245 -244 246 -243
rect 246 -244 247 -243
rect 247 -244 248 -243
rect 248 -244 249 -243
rect 249 -244 250 -243
rect 250 -244 251 -243
rect 251 -244 252 -243
rect 252 -244 253 -243
rect 253 -244 254 -243
rect 254 -244 255 -243
rect 255 -244 256 -243
rect 256 -244 257 -243
rect 257 -244 258 -243
rect 258 -244 259 -243
rect 259 -244 260 -243
rect 260 -244 261 -243
rect 261 -244 262 -243
rect 262 -244 263 -243
rect 263 -244 264 -243
rect 264 -244 265 -243
rect 265 -244 266 -243
rect 266 -244 267 -243
rect 267 -244 268 -243
rect 268 -244 269 -243
rect 269 -244 270 -243
rect 270 -244 271 -243
rect 271 -244 272 -243
rect 272 -244 273 -243
rect 273 -244 274 -243
rect 274 -244 275 -243
rect 275 -244 276 -243
rect 276 -244 277 -243
rect 277 -244 278 -243
rect 278 -244 279 -243
rect 279 -244 280 -243
rect 280 -244 281 -243
rect 281 -244 282 -243
rect 282 -244 283 -243
rect 283 -244 284 -243
rect 284 -244 285 -243
rect 285 -244 286 -243
rect 286 -244 287 -243
rect 287 -244 288 -243
rect 288 -244 289 -243
rect 289 -244 290 -243
rect 290 -244 291 -243
rect 291 -244 292 -243
rect 292 -244 293 -243
rect 293 -244 294 -243
rect 294 -244 295 -243
rect 295 -244 296 -243
rect 296 -244 297 -243
rect 297 -244 298 -243
rect 298 -244 299 -243
rect 299 -244 300 -243
rect 300 -244 301 -243
rect 301 -244 302 -243
rect 302 -244 303 -243
rect 303 -244 304 -243
rect 304 -244 305 -243
rect 305 -244 306 -243
rect 306 -244 307 -243
rect 307 -244 308 -243
rect 308 -244 309 -243
rect 309 -244 310 -243
rect 310 -244 311 -243
rect 311 -244 312 -243
rect 312 -244 313 -243
rect 313 -244 314 -243
rect 314 -244 315 -243
rect 315 -244 316 -243
rect 316 -244 317 -243
rect 317 -244 318 -243
rect 318 -244 319 -243
rect 319 -244 320 -243
rect 320 -244 321 -243
rect 321 -244 322 -243
rect 322 -244 323 -243
rect 323 -244 324 -243
rect 324 -244 325 -243
rect 325 -244 326 -243
rect 326 -244 327 -243
rect 327 -244 328 -243
rect 328 -244 329 -243
rect 329 -244 330 -243
rect 330 -244 331 -243
rect 331 -244 332 -243
rect 332 -244 333 -243
rect 333 -244 334 -243
rect 334 -244 335 -243
rect 335 -244 336 -243
rect 336 -244 337 -243
rect 337 -244 338 -243
rect 338 -244 339 -243
rect 339 -244 340 -243
rect 340 -244 341 -243
rect 341 -244 342 -243
rect 342 -244 343 -243
rect 343 -244 344 -243
rect 344 -244 345 -243
rect 345 -244 346 -243
rect 346 -244 347 -243
rect 347 -244 348 -243
rect 348 -244 349 -243
rect 349 -244 350 -243
rect 350 -244 351 -243
rect 351 -244 352 -243
rect 352 -244 353 -243
rect 353 -244 354 -243
rect 354 -244 355 -243
rect 355 -244 356 -243
rect 356 -244 357 -243
rect 357 -244 358 -243
rect 358 -244 359 -243
rect 359 -244 360 -243
rect 360 -244 361 -243
rect 361 -244 362 -243
rect 362 -244 363 -243
rect 363 -244 364 -243
rect 364 -244 365 -243
rect 365 -244 366 -243
rect 366 -244 367 -243
rect 367 -244 368 -243
rect 368 -244 369 -243
rect 369 -244 370 -243
rect 370 -244 371 -243
rect 371 -244 372 -243
rect 372 -244 373 -243
rect 373 -244 374 -243
rect 374 -244 375 -243
rect 375 -244 376 -243
rect 376 -244 377 -243
rect 377 -244 378 -243
rect 378 -244 379 -243
rect 379 -244 380 -243
rect 380 -244 381 -243
rect 381 -244 382 -243
rect 382 -244 383 -243
rect 383 -244 384 -243
rect 384 -244 385 -243
rect 385 -244 386 -243
rect 386 -244 387 -243
rect 387 -244 388 -243
rect 388 -244 389 -243
rect 389 -244 390 -243
rect 390 -244 391 -243
rect 391 -244 392 -243
rect 392 -244 393 -243
rect 393 -244 394 -243
rect 394 -244 395 -243
rect 395 -244 396 -243
rect 396 -244 397 -243
rect 397 -244 398 -243
rect 398 -244 399 -243
rect 399 -244 400 -243
rect 400 -244 401 -243
rect 401 -244 402 -243
rect 402 -244 403 -243
rect 403 -244 404 -243
rect 404 -244 405 -243
rect 405 -244 406 -243
rect 406 -244 407 -243
rect 407 -244 408 -243
rect 408 -244 409 -243
rect 409 -244 410 -243
rect 410 -244 411 -243
rect 411 -244 412 -243
rect 412 -244 413 -243
rect 413 -244 414 -243
rect 414 -244 415 -243
rect 415 -244 416 -243
rect 416 -244 417 -243
rect 417 -244 418 -243
rect 418 -244 419 -243
rect 419 -244 420 -243
rect 420 -244 421 -243
rect 421 -244 422 -243
rect 422 -244 423 -243
rect 423 -244 424 -243
rect 424 -244 425 -243
rect 425 -244 426 -243
rect 426 -244 427 -243
rect 427 -244 428 -243
rect 428 -244 429 -243
rect 429 -244 430 -243
rect 430 -244 431 -243
rect 431 -244 432 -243
rect 432 -244 433 -243
rect 433 -244 434 -243
rect 434 -244 435 -243
rect 435 -244 436 -243
rect 436 -244 437 -243
rect 437 -244 438 -243
rect 438 -244 439 -243
rect 439 -244 440 -243
rect 440 -244 441 -243
rect 441 -244 442 -243
rect 442 -244 443 -243
rect 443 -244 444 -243
rect 444 -244 445 -243
rect 445 -244 446 -243
rect 446 -244 447 -243
rect 447 -244 448 -243
rect 448 -244 449 -243
rect 449 -244 450 -243
rect 450 -244 451 -243
rect 451 -244 452 -243
rect 452 -244 453 -243
rect 453 -244 454 -243
rect 454 -244 455 -243
rect 455 -244 456 -243
rect 456 -244 457 -243
rect 457 -244 458 -243
rect 458 -244 459 -243
rect 459 -244 460 -243
rect 460 -244 461 -243
rect 461 -244 462 -243
rect 462 -244 463 -243
rect 463 -244 464 -243
rect 464 -244 465 -243
rect 465 -244 466 -243
rect 466 -244 467 -243
rect 467 -244 468 -243
rect 468 -244 469 -243
rect 469 -244 470 -243
rect 470 -244 471 -243
rect 471 -244 472 -243
rect 472 -244 473 -243
rect 473 -244 474 -243
rect 474 -244 475 -243
rect 475 -244 476 -243
rect 476 -244 477 -243
rect 477 -244 478 -243
rect 478 -244 479 -243
rect 479 -244 480 -243
rect 2 -245 3 -244
rect 3 -245 4 -244
rect 4 -245 5 -244
rect 5 -245 6 -244
rect 6 -245 7 -244
rect 7 -245 8 -244
rect 8 -245 9 -244
rect 9 -245 10 -244
rect 10 -245 11 -244
rect 11 -245 12 -244
rect 12 -245 13 -244
rect 13 -245 14 -244
rect 14 -245 15 -244
rect 15 -245 16 -244
rect 16 -245 17 -244
rect 17 -245 18 -244
rect 18 -245 19 -244
rect 19 -245 20 -244
rect 20 -245 21 -244
rect 21 -245 22 -244
rect 22 -245 23 -244
rect 23 -245 24 -244
rect 24 -245 25 -244
rect 25 -245 26 -244
rect 26 -245 27 -244
rect 27 -245 28 -244
rect 28 -245 29 -244
rect 29 -245 30 -244
rect 30 -245 31 -244
rect 31 -245 32 -244
rect 32 -245 33 -244
rect 33 -245 34 -244
rect 34 -245 35 -244
rect 35 -245 36 -244
rect 36 -245 37 -244
rect 37 -245 38 -244
rect 38 -245 39 -244
rect 39 -245 40 -244
rect 40 -245 41 -244
rect 41 -245 42 -244
rect 42 -245 43 -244
rect 43 -245 44 -244
rect 44 -245 45 -244
rect 45 -245 46 -244
rect 46 -245 47 -244
rect 47 -245 48 -244
rect 48 -245 49 -244
rect 49 -245 50 -244
rect 50 -245 51 -244
rect 51 -245 52 -244
rect 52 -245 53 -244
rect 53 -245 54 -244
rect 54 -245 55 -244
rect 55 -245 56 -244
rect 56 -245 57 -244
rect 57 -245 58 -244
rect 58 -245 59 -244
rect 59 -245 60 -244
rect 60 -245 61 -244
rect 61 -245 62 -244
rect 62 -245 63 -244
rect 63 -245 64 -244
rect 64 -245 65 -244
rect 65 -245 66 -244
rect 66 -245 67 -244
rect 67 -245 68 -244
rect 68 -245 69 -244
rect 69 -245 70 -244
rect 70 -245 71 -244
rect 71 -245 72 -244
rect 72 -245 73 -244
rect 73 -245 74 -244
rect 74 -245 75 -244
rect 75 -245 76 -244
rect 76 -245 77 -244
rect 77 -245 78 -244
rect 78 -245 79 -244
rect 79 -245 80 -244
rect 80 -245 81 -244
rect 81 -245 82 -244
rect 82 -245 83 -244
rect 83 -245 84 -244
rect 84 -245 85 -244
rect 85 -245 86 -244
rect 86 -245 87 -244
rect 87 -245 88 -244
rect 88 -245 89 -244
rect 89 -245 90 -244
rect 90 -245 91 -244
rect 91 -245 92 -244
rect 92 -245 93 -244
rect 93 -245 94 -244
rect 94 -245 95 -244
rect 95 -245 96 -244
rect 96 -245 97 -244
rect 97 -245 98 -244
rect 98 -245 99 -244
rect 99 -245 100 -244
rect 100 -245 101 -244
rect 101 -245 102 -244
rect 102 -245 103 -244
rect 103 -245 104 -244
rect 104 -245 105 -244
rect 105 -245 106 -244
rect 106 -245 107 -244
rect 107 -245 108 -244
rect 108 -245 109 -244
rect 109 -245 110 -244
rect 110 -245 111 -244
rect 111 -245 112 -244
rect 112 -245 113 -244
rect 113 -245 114 -244
rect 114 -245 115 -244
rect 115 -245 116 -244
rect 116 -245 117 -244
rect 117 -245 118 -244
rect 118 -245 119 -244
rect 119 -245 120 -244
rect 120 -245 121 -244
rect 121 -245 122 -244
rect 122 -245 123 -244
rect 123 -245 124 -244
rect 124 -245 125 -244
rect 125 -245 126 -244
rect 126 -245 127 -244
rect 127 -245 128 -244
rect 128 -245 129 -244
rect 129 -245 130 -244
rect 130 -245 131 -244
rect 131 -245 132 -244
rect 132 -245 133 -244
rect 133 -245 134 -244
rect 134 -245 135 -244
rect 135 -245 136 -244
rect 136 -245 137 -244
rect 137 -245 138 -244
rect 138 -245 139 -244
rect 139 -245 140 -244
rect 140 -245 141 -244
rect 141 -245 142 -244
rect 142 -245 143 -244
rect 143 -245 144 -244
rect 144 -245 145 -244
rect 145 -245 146 -244
rect 146 -245 147 -244
rect 147 -245 148 -244
rect 148 -245 149 -244
rect 149 -245 150 -244
rect 150 -245 151 -244
rect 151 -245 152 -244
rect 152 -245 153 -244
rect 153 -245 154 -244
rect 154 -245 155 -244
rect 155 -245 156 -244
rect 156 -245 157 -244
rect 157 -245 158 -244
rect 158 -245 159 -244
rect 159 -245 160 -244
rect 160 -245 161 -244
rect 161 -245 162 -244
rect 162 -245 163 -244
rect 163 -245 164 -244
rect 164 -245 165 -244
rect 165 -245 166 -244
rect 166 -245 167 -244
rect 167 -245 168 -244
rect 168 -245 169 -244
rect 169 -245 170 -244
rect 170 -245 171 -244
rect 171 -245 172 -244
rect 172 -245 173 -244
rect 173 -245 174 -244
rect 174 -245 175 -244
rect 175 -245 176 -244
rect 176 -245 177 -244
rect 177 -245 178 -244
rect 178 -245 179 -244
rect 179 -245 180 -244
rect 180 -245 181 -244
rect 181 -245 182 -244
rect 182 -245 183 -244
rect 183 -245 184 -244
rect 184 -245 185 -244
rect 185 -245 186 -244
rect 186 -245 187 -244
rect 187 -245 188 -244
rect 188 -245 189 -244
rect 189 -245 190 -244
rect 190 -245 191 -244
rect 191 -245 192 -244
rect 192 -245 193 -244
rect 193 -245 194 -244
rect 194 -245 195 -244
rect 195 -245 196 -244
rect 196 -245 197 -244
rect 197 -245 198 -244
rect 198 -245 199 -244
rect 199 -245 200 -244
rect 200 -245 201 -244
rect 201 -245 202 -244
rect 202 -245 203 -244
rect 203 -245 204 -244
rect 204 -245 205 -244
rect 205 -245 206 -244
rect 206 -245 207 -244
rect 207 -245 208 -244
rect 208 -245 209 -244
rect 209 -245 210 -244
rect 210 -245 211 -244
rect 211 -245 212 -244
rect 212 -245 213 -244
rect 213 -245 214 -244
rect 214 -245 215 -244
rect 215 -245 216 -244
rect 216 -245 217 -244
rect 217 -245 218 -244
rect 218 -245 219 -244
rect 219 -245 220 -244
rect 220 -245 221 -244
rect 221 -245 222 -244
rect 222 -245 223 -244
rect 223 -245 224 -244
rect 224 -245 225 -244
rect 225 -245 226 -244
rect 226 -245 227 -244
rect 227 -245 228 -244
rect 228 -245 229 -244
rect 229 -245 230 -244
rect 230 -245 231 -244
rect 231 -245 232 -244
rect 232 -245 233 -244
rect 233 -245 234 -244
rect 234 -245 235 -244
rect 235 -245 236 -244
rect 236 -245 237 -244
rect 237 -245 238 -244
rect 238 -245 239 -244
rect 239 -245 240 -244
rect 240 -245 241 -244
rect 241 -245 242 -244
rect 242 -245 243 -244
rect 243 -245 244 -244
rect 244 -245 245 -244
rect 245 -245 246 -244
rect 246 -245 247 -244
rect 247 -245 248 -244
rect 248 -245 249 -244
rect 249 -245 250 -244
rect 250 -245 251 -244
rect 251 -245 252 -244
rect 252 -245 253 -244
rect 253 -245 254 -244
rect 254 -245 255 -244
rect 255 -245 256 -244
rect 256 -245 257 -244
rect 257 -245 258 -244
rect 258 -245 259 -244
rect 259 -245 260 -244
rect 260 -245 261 -244
rect 261 -245 262 -244
rect 262 -245 263 -244
rect 263 -245 264 -244
rect 264 -245 265 -244
rect 265 -245 266 -244
rect 266 -245 267 -244
rect 267 -245 268 -244
rect 268 -245 269 -244
rect 269 -245 270 -244
rect 270 -245 271 -244
rect 271 -245 272 -244
rect 272 -245 273 -244
rect 273 -245 274 -244
rect 274 -245 275 -244
rect 275 -245 276 -244
rect 276 -245 277 -244
rect 277 -245 278 -244
rect 278 -245 279 -244
rect 279 -245 280 -244
rect 280 -245 281 -244
rect 281 -245 282 -244
rect 282 -245 283 -244
rect 283 -245 284 -244
rect 284 -245 285 -244
rect 285 -245 286 -244
rect 286 -245 287 -244
rect 287 -245 288 -244
rect 288 -245 289 -244
rect 289 -245 290 -244
rect 290 -245 291 -244
rect 291 -245 292 -244
rect 292 -245 293 -244
rect 293 -245 294 -244
rect 294 -245 295 -244
rect 295 -245 296 -244
rect 296 -245 297 -244
rect 297 -245 298 -244
rect 298 -245 299 -244
rect 299 -245 300 -244
rect 300 -245 301 -244
rect 301 -245 302 -244
rect 302 -245 303 -244
rect 303 -245 304 -244
rect 304 -245 305 -244
rect 305 -245 306 -244
rect 306 -245 307 -244
rect 307 -245 308 -244
rect 308 -245 309 -244
rect 309 -245 310 -244
rect 310 -245 311 -244
rect 311 -245 312 -244
rect 312 -245 313 -244
rect 313 -245 314 -244
rect 314 -245 315 -244
rect 315 -245 316 -244
rect 316 -245 317 -244
rect 317 -245 318 -244
rect 318 -245 319 -244
rect 319 -245 320 -244
rect 320 -245 321 -244
rect 321 -245 322 -244
rect 322 -245 323 -244
rect 323 -245 324 -244
rect 324 -245 325 -244
rect 325 -245 326 -244
rect 326 -245 327 -244
rect 327 -245 328 -244
rect 328 -245 329 -244
rect 329 -245 330 -244
rect 330 -245 331 -244
rect 331 -245 332 -244
rect 332 -245 333 -244
rect 333 -245 334 -244
rect 334 -245 335 -244
rect 335 -245 336 -244
rect 336 -245 337 -244
rect 337 -245 338 -244
rect 338 -245 339 -244
rect 339 -245 340 -244
rect 340 -245 341 -244
rect 341 -245 342 -244
rect 342 -245 343 -244
rect 343 -245 344 -244
rect 344 -245 345 -244
rect 345 -245 346 -244
rect 346 -245 347 -244
rect 347 -245 348 -244
rect 348 -245 349 -244
rect 349 -245 350 -244
rect 350 -245 351 -244
rect 351 -245 352 -244
rect 352 -245 353 -244
rect 353 -245 354 -244
rect 354 -245 355 -244
rect 355 -245 356 -244
rect 356 -245 357 -244
rect 357 -245 358 -244
rect 358 -245 359 -244
rect 359 -245 360 -244
rect 360 -245 361 -244
rect 361 -245 362 -244
rect 362 -245 363 -244
rect 363 -245 364 -244
rect 364 -245 365 -244
rect 365 -245 366 -244
rect 366 -245 367 -244
rect 367 -245 368 -244
rect 368 -245 369 -244
rect 369 -245 370 -244
rect 370 -245 371 -244
rect 371 -245 372 -244
rect 372 -245 373 -244
rect 373 -245 374 -244
rect 374 -245 375 -244
rect 375 -245 376 -244
rect 376 -245 377 -244
rect 377 -245 378 -244
rect 378 -245 379 -244
rect 379 -245 380 -244
rect 380 -245 381 -244
rect 381 -245 382 -244
rect 382 -245 383 -244
rect 383 -245 384 -244
rect 384 -245 385 -244
rect 385 -245 386 -244
rect 386 -245 387 -244
rect 387 -245 388 -244
rect 388 -245 389 -244
rect 389 -245 390 -244
rect 390 -245 391 -244
rect 391 -245 392 -244
rect 392 -245 393 -244
rect 393 -245 394 -244
rect 394 -245 395 -244
rect 395 -245 396 -244
rect 396 -245 397 -244
rect 397 -245 398 -244
rect 398 -245 399 -244
rect 399 -245 400 -244
rect 400 -245 401 -244
rect 401 -245 402 -244
rect 402 -245 403 -244
rect 403 -245 404 -244
rect 404 -245 405 -244
rect 405 -245 406 -244
rect 406 -245 407 -244
rect 407 -245 408 -244
rect 408 -245 409 -244
rect 409 -245 410 -244
rect 410 -245 411 -244
rect 411 -245 412 -244
rect 412 -245 413 -244
rect 413 -245 414 -244
rect 414 -245 415 -244
rect 415 -245 416 -244
rect 416 -245 417 -244
rect 417 -245 418 -244
rect 418 -245 419 -244
rect 419 -245 420 -244
rect 420 -245 421 -244
rect 421 -245 422 -244
rect 422 -245 423 -244
rect 423 -245 424 -244
rect 424 -245 425 -244
rect 425 -245 426 -244
rect 426 -245 427 -244
rect 427 -245 428 -244
rect 428 -245 429 -244
rect 429 -245 430 -244
rect 430 -245 431 -244
rect 431 -245 432 -244
rect 432 -245 433 -244
rect 433 -245 434 -244
rect 434 -245 435 -244
rect 435 -245 436 -244
rect 436 -245 437 -244
rect 437 -245 438 -244
rect 438 -245 439 -244
rect 439 -245 440 -244
rect 440 -245 441 -244
rect 441 -245 442 -244
rect 442 -245 443 -244
rect 443 -245 444 -244
rect 444 -245 445 -244
rect 445 -245 446 -244
rect 446 -245 447 -244
rect 447 -245 448 -244
rect 448 -245 449 -244
rect 449 -245 450 -244
rect 450 -245 451 -244
rect 451 -245 452 -244
rect 452 -245 453 -244
rect 453 -245 454 -244
rect 454 -245 455 -244
rect 455 -245 456 -244
rect 456 -245 457 -244
rect 457 -245 458 -244
rect 458 -245 459 -244
rect 459 -245 460 -244
rect 460 -245 461 -244
rect 461 -245 462 -244
rect 462 -245 463 -244
rect 463 -245 464 -244
rect 464 -245 465 -244
rect 465 -245 466 -244
rect 466 -245 467 -244
rect 467 -245 468 -244
rect 468 -245 469 -244
rect 469 -245 470 -244
rect 470 -245 471 -244
rect 471 -245 472 -244
rect 472 -245 473 -244
rect 473 -245 474 -244
rect 474 -245 475 -244
rect 475 -245 476 -244
rect 476 -245 477 -244
rect 477 -245 478 -244
rect 478 -245 479 -244
rect 479 -245 480 -244
rect 2 -246 3 -245
rect 3 -246 4 -245
rect 4 -246 5 -245
rect 5 -246 6 -245
rect 6 -246 7 -245
rect 7 -246 8 -245
rect 8 -246 9 -245
rect 9 -246 10 -245
rect 10 -246 11 -245
rect 11 -246 12 -245
rect 12 -246 13 -245
rect 13 -246 14 -245
rect 14 -246 15 -245
rect 15 -246 16 -245
rect 16 -246 17 -245
rect 17 -246 18 -245
rect 18 -246 19 -245
rect 19 -246 20 -245
rect 20 -246 21 -245
rect 21 -246 22 -245
rect 22 -246 23 -245
rect 23 -246 24 -245
rect 24 -246 25 -245
rect 25 -246 26 -245
rect 26 -246 27 -245
rect 27 -246 28 -245
rect 28 -246 29 -245
rect 29 -246 30 -245
rect 30 -246 31 -245
rect 31 -246 32 -245
rect 32 -246 33 -245
rect 33 -246 34 -245
rect 34 -246 35 -245
rect 35 -246 36 -245
rect 36 -246 37 -245
rect 37 -246 38 -245
rect 38 -246 39 -245
rect 39 -246 40 -245
rect 40 -246 41 -245
rect 41 -246 42 -245
rect 42 -246 43 -245
rect 43 -246 44 -245
rect 44 -246 45 -245
rect 45 -246 46 -245
rect 46 -246 47 -245
rect 47 -246 48 -245
rect 48 -246 49 -245
rect 49 -246 50 -245
rect 50 -246 51 -245
rect 51 -246 52 -245
rect 52 -246 53 -245
rect 53 -246 54 -245
rect 54 -246 55 -245
rect 55 -246 56 -245
rect 56 -246 57 -245
rect 57 -246 58 -245
rect 58 -246 59 -245
rect 59 -246 60 -245
rect 60 -246 61 -245
rect 61 -246 62 -245
rect 62 -246 63 -245
rect 63 -246 64 -245
rect 64 -246 65 -245
rect 65 -246 66 -245
rect 66 -246 67 -245
rect 67 -246 68 -245
rect 68 -246 69 -245
rect 69 -246 70 -245
rect 70 -246 71 -245
rect 71 -246 72 -245
rect 72 -246 73 -245
rect 73 -246 74 -245
rect 74 -246 75 -245
rect 75 -246 76 -245
rect 76 -246 77 -245
rect 77 -246 78 -245
rect 78 -246 79 -245
rect 79 -246 80 -245
rect 80 -246 81 -245
rect 81 -246 82 -245
rect 82 -246 83 -245
rect 83 -246 84 -245
rect 84 -246 85 -245
rect 85 -246 86 -245
rect 86 -246 87 -245
rect 87 -246 88 -245
rect 88 -246 89 -245
rect 89 -246 90 -245
rect 90 -246 91 -245
rect 91 -246 92 -245
rect 92 -246 93 -245
rect 93 -246 94 -245
rect 94 -246 95 -245
rect 95 -246 96 -245
rect 96 -246 97 -245
rect 97 -246 98 -245
rect 98 -246 99 -245
rect 99 -246 100 -245
rect 100 -246 101 -245
rect 101 -246 102 -245
rect 102 -246 103 -245
rect 103 -246 104 -245
rect 104 -246 105 -245
rect 105 -246 106 -245
rect 106 -246 107 -245
rect 107 -246 108 -245
rect 108 -246 109 -245
rect 109 -246 110 -245
rect 110 -246 111 -245
rect 111 -246 112 -245
rect 112 -246 113 -245
rect 113 -246 114 -245
rect 114 -246 115 -245
rect 115 -246 116 -245
rect 116 -246 117 -245
rect 117 -246 118 -245
rect 118 -246 119 -245
rect 119 -246 120 -245
rect 120 -246 121 -245
rect 121 -246 122 -245
rect 122 -246 123 -245
rect 123 -246 124 -245
rect 124 -246 125 -245
rect 125 -246 126 -245
rect 126 -246 127 -245
rect 127 -246 128 -245
rect 128 -246 129 -245
rect 129 -246 130 -245
rect 130 -246 131 -245
rect 131 -246 132 -245
rect 132 -246 133 -245
rect 133 -246 134 -245
rect 134 -246 135 -245
rect 135 -246 136 -245
rect 136 -246 137 -245
rect 137 -246 138 -245
rect 138 -246 139 -245
rect 139 -246 140 -245
rect 140 -246 141 -245
rect 141 -246 142 -245
rect 142 -246 143 -245
rect 143 -246 144 -245
rect 144 -246 145 -245
rect 145 -246 146 -245
rect 146 -246 147 -245
rect 147 -246 148 -245
rect 148 -246 149 -245
rect 149 -246 150 -245
rect 150 -246 151 -245
rect 151 -246 152 -245
rect 152 -246 153 -245
rect 153 -246 154 -245
rect 154 -246 155 -245
rect 155 -246 156 -245
rect 156 -246 157 -245
rect 157 -246 158 -245
rect 158 -246 159 -245
rect 159 -246 160 -245
rect 160 -246 161 -245
rect 161 -246 162 -245
rect 162 -246 163 -245
rect 163 -246 164 -245
rect 164 -246 165 -245
rect 165 -246 166 -245
rect 166 -246 167 -245
rect 167 -246 168 -245
rect 168 -246 169 -245
rect 169 -246 170 -245
rect 170 -246 171 -245
rect 171 -246 172 -245
rect 172 -246 173 -245
rect 173 -246 174 -245
rect 174 -246 175 -245
rect 175 -246 176 -245
rect 176 -246 177 -245
rect 177 -246 178 -245
rect 178 -246 179 -245
rect 179 -246 180 -245
rect 180 -246 181 -245
rect 181 -246 182 -245
rect 182 -246 183 -245
rect 183 -246 184 -245
rect 184 -246 185 -245
rect 185 -246 186 -245
rect 186 -246 187 -245
rect 187 -246 188 -245
rect 188 -246 189 -245
rect 189 -246 190 -245
rect 190 -246 191 -245
rect 191 -246 192 -245
rect 192 -246 193 -245
rect 193 -246 194 -245
rect 194 -246 195 -245
rect 195 -246 196 -245
rect 196 -246 197 -245
rect 197 -246 198 -245
rect 198 -246 199 -245
rect 199 -246 200 -245
rect 200 -246 201 -245
rect 201 -246 202 -245
rect 202 -246 203 -245
rect 203 -246 204 -245
rect 204 -246 205 -245
rect 205 -246 206 -245
rect 206 -246 207 -245
rect 207 -246 208 -245
rect 208 -246 209 -245
rect 209 -246 210 -245
rect 210 -246 211 -245
rect 211 -246 212 -245
rect 212 -246 213 -245
rect 213 -246 214 -245
rect 214 -246 215 -245
rect 215 -246 216 -245
rect 216 -246 217 -245
rect 217 -246 218 -245
rect 218 -246 219 -245
rect 219 -246 220 -245
rect 220 -246 221 -245
rect 221 -246 222 -245
rect 222 -246 223 -245
rect 223 -246 224 -245
rect 224 -246 225 -245
rect 225 -246 226 -245
rect 226 -246 227 -245
rect 227 -246 228 -245
rect 228 -246 229 -245
rect 229 -246 230 -245
rect 230 -246 231 -245
rect 231 -246 232 -245
rect 232 -246 233 -245
rect 233 -246 234 -245
rect 234 -246 235 -245
rect 235 -246 236 -245
rect 236 -246 237 -245
rect 237 -246 238 -245
rect 238 -246 239 -245
rect 239 -246 240 -245
rect 240 -246 241 -245
rect 241 -246 242 -245
rect 242 -246 243 -245
rect 243 -246 244 -245
rect 244 -246 245 -245
rect 245 -246 246 -245
rect 246 -246 247 -245
rect 247 -246 248 -245
rect 248 -246 249 -245
rect 249 -246 250 -245
rect 250 -246 251 -245
rect 251 -246 252 -245
rect 252 -246 253 -245
rect 253 -246 254 -245
rect 254 -246 255 -245
rect 255 -246 256 -245
rect 256 -246 257 -245
rect 257 -246 258 -245
rect 258 -246 259 -245
rect 259 -246 260 -245
rect 260 -246 261 -245
rect 261 -246 262 -245
rect 262 -246 263 -245
rect 263 -246 264 -245
rect 264 -246 265 -245
rect 265 -246 266 -245
rect 266 -246 267 -245
rect 267 -246 268 -245
rect 268 -246 269 -245
rect 269 -246 270 -245
rect 270 -246 271 -245
rect 271 -246 272 -245
rect 272 -246 273 -245
rect 273 -246 274 -245
rect 274 -246 275 -245
rect 275 -246 276 -245
rect 276 -246 277 -245
rect 277 -246 278 -245
rect 278 -246 279 -245
rect 279 -246 280 -245
rect 280 -246 281 -245
rect 281 -246 282 -245
rect 282 -246 283 -245
rect 283 -246 284 -245
rect 284 -246 285 -245
rect 285 -246 286 -245
rect 286 -246 287 -245
rect 287 -246 288 -245
rect 288 -246 289 -245
rect 289 -246 290 -245
rect 290 -246 291 -245
rect 291 -246 292 -245
rect 292 -246 293 -245
rect 293 -246 294 -245
rect 294 -246 295 -245
rect 295 -246 296 -245
rect 296 -246 297 -245
rect 297 -246 298 -245
rect 298 -246 299 -245
rect 299 -246 300 -245
rect 300 -246 301 -245
rect 301 -246 302 -245
rect 302 -246 303 -245
rect 303 -246 304 -245
rect 304 -246 305 -245
rect 305 -246 306 -245
rect 306 -246 307 -245
rect 307 -246 308 -245
rect 308 -246 309 -245
rect 309 -246 310 -245
rect 310 -246 311 -245
rect 311 -246 312 -245
rect 312 -246 313 -245
rect 313 -246 314 -245
rect 314 -246 315 -245
rect 315 -246 316 -245
rect 316 -246 317 -245
rect 317 -246 318 -245
rect 318 -246 319 -245
rect 319 -246 320 -245
rect 320 -246 321 -245
rect 321 -246 322 -245
rect 322 -246 323 -245
rect 323 -246 324 -245
rect 324 -246 325 -245
rect 325 -246 326 -245
rect 326 -246 327 -245
rect 327 -246 328 -245
rect 328 -246 329 -245
rect 329 -246 330 -245
rect 330 -246 331 -245
rect 331 -246 332 -245
rect 332 -246 333 -245
rect 333 -246 334 -245
rect 334 -246 335 -245
rect 335 -246 336 -245
rect 336 -246 337 -245
rect 337 -246 338 -245
rect 338 -246 339 -245
rect 339 -246 340 -245
rect 340 -246 341 -245
rect 341 -246 342 -245
rect 342 -246 343 -245
rect 343 -246 344 -245
rect 344 -246 345 -245
rect 345 -246 346 -245
rect 346 -246 347 -245
rect 347 -246 348 -245
rect 348 -246 349 -245
rect 349 -246 350 -245
rect 350 -246 351 -245
rect 351 -246 352 -245
rect 352 -246 353 -245
rect 353 -246 354 -245
rect 354 -246 355 -245
rect 355 -246 356 -245
rect 356 -246 357 -245
rect 357 -246 358 -245
rect 358 -246 359 -245
rect 359 -246 360 -245
rect 360 -246 361 -245
rect 361 -246 362 -245
rect 362 -246 363 -245
rect 363 -246 364 -245
rect 364 -246 365 -245
rect 365 -246 366 -245
rect 366 -246 367 -245
rect 367 -246 368 -245
rect 368 -246 369 -245
rect 369 -246 370 -245
rect 370 -246 371 -245
rect 371 -246 372 -245
rect 372 -246 373 -245
rect 373 -246 374 -245
rect 374 -246 375 -245
rect 375 -246 376 -245
rect 376 -246 377 -245
rect 377 -246 378 -245
rect 378 -246 379 -245
rect 379 -246 380 -245
rect 380 -246 381 -245
rect 381 -246 382 -245
rect 382 -246 383 -245
rect 383 -246 384 -245
rect 384 -246 385 -245
rect 385 -246 386 -245
rect 386 -246 387 -245
rect 387 -246 388 -245
rect 388 -246 389 -245
rect 389 -246 390 -245
rect 390 -246 391 -245
rect 391 -246 392 -245
rect 392 -246 393 -245
rect 393 -246 394 -245
rect 394 -246 395 -245
rect 395 -246 396 -245
rect 396 -246 397 -245
rect 397 -246 398 -245
rect 398 -246 399 -245
rect 399 -246 400 -245
rect 400 -246 401 -245
rect 401 -246 402 -245
rect 402 -246 403 -245
rect 403 -246 404 -245
rect 404 -246 405 -245
rect 405 -246 406 -245
rect 406 -246 407 -245
rect 407 -246 408 -245
rect 408 -246 409 -245
rect 409 -246 410 -245
rect 410 -246 411 -245
rect 411 -246 412 -245
rect 412 -246 413 -245
rect 413 -246 414 -245
rect 414 -246 415 -245
rect 415 -246 416 -245
rect 416 -246 417 -245
rect 417 -246 418 -245
rect 418 -246 419 -245
rect 419 -246 420 -245
rect 420 -246 421 -245
rect 421 -246 422 -245
rect 422 -246 423 -245
rect 423 -246 424 -245
rect 424 -246 425 -245
rect 425 -246 426 -245
rect 426 -246 427 -245
rect 427 -246 428 -245
rect 428 -246 429 -245
rect 429 -246 430 -245
rect 430 -246 431 -245
rect 431 -246 432 -245
rect 432 -246 433 -245
rect 433 -246 434 -245
rect 434 -246 435 -245
rect 435 -246 436 -245
rect 436 -246 437 -245
rect 437 -246 438 -245
rect 438 -246 439 -245
rect 439 -246 440 -245
rect 440 -246 441 -245
rect 441 -246 442 -245
rect 442 -246 443 -245
rect 443 -246 444 -245
rect 444 -246 445 -245
rect 445 -246 446 -245
rect 446 -246 447 -245
rect 447 -246 448 -245
rect 448 -246 449 -245
rect 449 -246 450 -245
rect 450 -246 451 -245
rect 451 -246 452 -245
rect 452 -246 453 -245
rect 453 -246 454 -245
rect 454 -246 455 -245
rect 455 -246 456 -245
rect 456 -246 457 -245
rect 457 -246 458 -245
rect 458 -246 459 -245
rect 459 -246 460 -245
rect 460 -246 461 -245
rect 461 -246 462 -245
rect 462 -246 463 -245
rect 463 -246 464 -245
rect 464 -246 465 -245
rect 465 -246 466 -245
rect 466 -246 467 -245
rect 467 -246 468 -245
rect 468 -246 469 -245
rect 469 -246 470 -245
rect 470 -246 471 -245
rect 471 -246 472 -245
rect 472 -246 473 -245
rect 473 -246 474 -245
rect 474 -246 475 -245
rect 475 -246 476 -245
rect 476 -246 477 -245
rect 477 -246 478 -245
rect 478 -246 479 -245
rect 479 -246 480 -245
rect 2 -247 3 -246
rect 3 -247 4 -246
rect 4 -247 5 -246
rect 5 -247 6 -246
rect 6 -247 7 -246
rect 7 -247 8 -246
rect 8 -247 9 -246
rect 9 -247 10 -246
rect 10 -247 11 -246
rect 11 -247 12 -246
rect 12 -247 13 -246
rect 13 -247 14 -246
rect 14 -247 15 -246
rect 15 -247 16 -246
rect 16 -247 17 -246
rect 17 -247 18 -246
rect 18 -247 19 -246
rect 19 -247 20 -246
rect 20 -247 21 -246
rect 21 -247 22 -246
rect 22 -247 23 -246
rect 23 -247 24 -246
rect 24 -247 25 -246
rect 25 -247 26 -246
rect 26 -247 27 -246
rect 27 -247 28 -246
rect 28 -247 29 -246
rect 29 -247 30 -246
rect 30 -247 31 -246
rect 31 -247 32 -246
rect 32 -247 33 -246
rect 33 -247 34 -246
rect 34 -247 35 -246
rect 35 -247 36 -246
rect 36 -247 37 -246
rect 37 -247 38 -246
rect 38 -247 39 -246
rect 39 -247 40 -246
rect 40 -247 41 -246
rect 41 -247 42 -246
rect 42 -247 43 -246
rect 43 -247 44 -246
rect 44 -247 45 -246
rect 45 -247 46 -246
rect 46 -247 47 -246
rect 47 -247 48 -246
rect 48 -247 49 -246
rect 49 -247 50 -246
rect 50 -247 51 -246
rect 51 -247 52 -246
rect 52 -247 53 -246
rect 53 -247 54 -246
rect 54 -247 55 -246
rect 55 -247 56 -246
rect 56 -247 57 -246
rect 57 -247 58 -246
rect 58 -247 59 -246
rect 59 -247 60 -246
rect 60 -247 61 -246
rect 61 -247 62 -246
rect 62 -247 63 -246
rect 63 -247 64 -246
rect 64 -247 65 -246
rect 65 -247 66 -246
rect 66 -247 67 -246
rect 67 -247 68 -246
rect 68 -247 69 -246
rect 69 -247 70 -246
rect 70 -247 71 -246
rect 71 -247 72 -246
rect 72 -247 73 -246
rect 73 -247 74 -246
rect 74 -247 75 -246
rect 75 -247 76 -246
rect 76 -247 77 -246
rect 77 -247 78 -246
rect 78 -247 79 -246
rect 79 -247 80 -246
rect 80 -247 81 -246
rect 81 -247 82 -246
rect 82 -247 83 -246
rect 83 -247 84 -246
rect 84 -247 85 -246
rect 85 -247 86 -246
rect 86 -247 87 -246
rect 87 -247 88 -246
rect 88 -247 89 -246
rect 89 -247 90 -246
rect 90 -247 91 -246
rect 91 -247 92 -246
rect 92 -247 93 -246
rect 93 -247 94 -246
rect 94 -247 95 -246
rect 95 -247 96 -246
rect 96 -247 97 -246
rect 97 -247 98 -246
rect 98 -247 99 -246
rect 99 -247 100 -246
rect 100 -247 101 -246
rect 101 -247 102 -246
rect 102 -247 103 -246
rect 103 -247 104 -246
rect 104 -247 105 -246
rect 105 -247 106 -246
rect 106 -247 107 -246
rect 107 -247 108 -246
rect 108 -247 109 -246
rect 109 -247 110 -246
rect 110 -247 111 -246
rect 111 -247 112 -246
rect 112 -247 113 -246
rect 113 -247 114 -246
rect 114 -247 115 -246
rect 115 -247 116 -246
rect 116 -247 117 -246
rect 117 -247 118 -246
rect 118 -247 119 -246
rect 119 -247 120 -246
rect 120 -247 121 -246
rect 121 -247 122 -246
rect 122 -247 123 -246
rect 123 -247 124 -246
rect 124 -247 125 -246
rect 125 -247 126 -246
rect 126 -247 127 -246
rect 127 -247 128 -246
rect 128 -247 129 -246
rect 129 -247 130 -246
rect 130 -247 131 -246
rect 131 -247 132 -246
rect 132 -247 133 -246
rect 133 -247 134 -246
rect 134 -247 135 -246
rect 135 -247 136 -246
rect 136 -247 137 -246
rect 137 -247 138 -246
rect 138 -247 139 -246
rect 139 -247 140 -246
rect 140 -247 141 -246
rect 141 -247 142 -246
rect 142 -247 143 -246
rect 143 -247 144 -246
rect 144 -247 145 -246
rect 145 -247 146 -246
rect 146 -247 147 -246
rect 147 -247 148 -246
rect 148 -247 149 -246
rect 149 -247 150 -246
rect 150 -247 151 -246
rect 151 -247 152 -246
rect 152 -247 153 -246
rect 153 -247 154 -246
rect 154 -247 155 -246
rect 155 -247 156 -246
rect 156 -247 157 -246
rect 157 -247 158 -246
rect 158 -247 159 -246
rect 159 -247 160 -246
rect 160 -247 161 -246
rect 161 -247 162 -246
rect 162 -247 163 -246
rect 163 -247 164 -246
rect 164 -247 165 -246
rect 165 -247 166 -246
rect 166 -247 167 -246
rect 167 -247 168 -246
rect 168 -247 169 -246
rect 169 -247 170 -246
rect 170 -247 171 -246
rect 171 -247 172 -246
rect 172 -247 173 -246
rect 173 -247 174 -246
rect 174 -247 175 -246
rect 175 -247 176 -246
rect 176 -247 177 -246
rect 177 -247 178 -246
rect 178 -247 179 -246
rect 179 -247 180 -246
rect 180 -247 181 -246
rect 181 -247 182 -246
rect 182 -247 183 -246
rect 183 -247 184 -246
rect 184 -247 185 -246
rect 185 -247 186 -246
rect 186 -247 187 -246
rect 187 -247 188 -246
rect 188 -247 189 -246
rect 189 -247 190 -246
rect 190 -247 191 -246
rect 191 -247 192 -246
rect 192 -247 193 -246
rect 193 -247 194 -246
rect 194 -247 195 -246
rect 195 -247 196 -246
rect 196 -247 197 -246
rect 197 -247 198 -246
rect 198 -247 199 -246
rect 199 -247 200 -246
rect 200 -247 201 -246
rect 201 -247 202 -246
rect 202 -247 203 -246
rect 203 -247 204 -246
rect 204 -247 205 -246
rect 205 -247 206 -246
rect 206 -247 207 -246
rect 207 -247 208 -246
rect 208 -247 209 -246
rect 209 -247 210 -246
rect 210 -247 211 -246
rect 211 -247 212 -246
rect 212 -247 213 -246
rect 213 -247 214 -246
rect 214 -247 215 -246
rect 215 -247 216 -246
rect 216 -247 217 -246
rect 217 -247 218 -246
rect 218 -247 219 -246
rect 219 -247 220 -246
rect 220 -247 221 -246
rect 221 -247 222 -246
rect 222 -247 223 -246
rect 223 -247 224 -246
rect 224 -247 225 -246
rect 225 -247 226 -246
rect 226 -247 227 -246
rect 227 -247 228 -246
rect 228 -247 229 -246
rect 229 -247 230 -246
rect 230 -247 231 -246
rect 231 -247 232 -246
rect 232 -247 233 -246
rect 233 -247 234 -246
rect 234 -247 235 -246
rect 235 -247 236 -246
rect 236 -247 237 -246
rect 237 -247 238 -246
rect 238 -247 239 -246
rect 239 -247 240 -246
rect 240 -247 241 -246
rect 241 -247 242 -246
rect 242 -247 243 -246
rect 243 -247 244 -246
rect 244 -247 245 -246
rect 245 -247 246 -246
rect 246 -247 247 -246
rect 247 -247 248 -246
rect 248 -247 249 -246
rect 249 -247 250 -246
rect 250 -247 251 -246
rect 251 -247 252 -246
rect 252 -247 253 -246
rect 253 -247 254 -246
rect 254 -247 255 -246
rect 255 -247 256 -246
rect 256 -247 257 -246
rect 257 -247 258 -246
rect 258 -247 259 -246
rect 259 -247 260 -246
rect 260 -247 261 -246
rect 261 -247 262 -246
rect 262 -247 263 -246
rect 263 -247 264 -246
rect 264 -247 265 -246
rect 265 -247 266 -246
rect 266 -247 267 -246
rect 267 -247 268 -246
rect 268 -247 269 -246
rect 269 -247 270 -246
rect 270 -247 271 -246
rect 271 -247 272 -246
rect 272 -247 273 -246
rect 273 -247 274 -246
rect 274 -247 275 -246
rect 275 -247 276 -246
rect 276 -247 277 -246
rect 277 -247 278 -246
rect 278 -247 279 -246
rect 279 -247 280 -246
rect 280 -247 281 -246
rect 281 -247 282 -246
rect 282 -247 283 -246
rect 283 -247 284 -246
rect 284 -247 285 -246
rect 285 -247 286 -246
rect 286 -247 287 -246
rect 287 -247 288 -246
rect 288 -247 289 -246
rect 289 -247 290 -246
rect 290 -247 291 -246
rect 291 -247 292 -246
rect 292 -247 293 -246
rect 293 -247 294 -246
rect 294 -247 295 -246
rect 295 -247 296 -246
rect 296 -247 297 -246
rect 297 -247 298 -246
rect 298 -247 299 -246
rect 299 -247 300 -246
rect 300 -247 301 -246
rect 301 -247 302 -246
rect 302 -247 303 -246
rect 303 -247 304 -246
rect 304 -247 305 -246
rect 305 -247 306 -246
rect 306 -247 307 -246
rect 307 -247 308 -246
rect 308 -247 309 -246
rect 309 -247 310 -246
rect 310 -247 311 -246
rect 311 -247 312 -246
rect 312 -247 313 -246
rect 313 -247 314 -246
rect 314 -247 315 -246
rect 315 -247 316 -246
rect 316 -247 317 -246
rect 317 -247 318 -246
rect 318 -247 319 -246
rect 319 -247 320 -246
rect 320 -247 321 -246
rect 321 -247 322 -246
rect 322 -247 323 -246
rect 323 -247 324 -246
rect 324 -247 325 -246
rect 325 -247 326 -246
rect 326 -247 327 -246
rect 327 -247 328 -246
rect 328 -247 329 -246
rect 329 -247 330 -246
rect 330 -247 331 -246
rect 331 -247 332 -246
rect 332 -247 333 -246
rect 333 -247 334 -246
rect 334 -247 335 -246
rect 335 -247 336 -246
rect 336 -247 337 -246
rect 337 -247 338 -246
rect 338 -247 339 -246
rect 339 -247 340 -246
rect 340 -247 341 -246
rect 341 -247 342 -246
rect 342 -247 343 -246
rect 343 -247 344 -246
rect 344 -247 345 -246
rect 345 -247 346 -246
rect 346 -247 347 -246
rect 347 -247 348 -246
rect 348 -247 349 -246
rect 349 -247 350 -246
rect 350 -247 351 -246
rect 351 -247 352 -246
rect 352 -247 353 -246
rect 353 -247 354 -246
rect 354 -247 355 -246
rect 355 -247 356 -246
rect 356 -247 357 -246
rect 357 -247 358 -246
rect 358 -247 359 -246
rect 359 -247 360 -246
rect 360 -247 361 -246
rect 361 -247 362 -246
rect 362 -247 363 -246
rect 363 -247 364 -246
rect 364 -247 365 -246
rect 365 -247 366 -246
rect 366 -247 367 -246
rect 367 -247 368 -246
rect 368 -247 369 -246
rect 369 -247 370 -246
rect 370 -247 371 -246
rect 371 -247 372 -246
rect 372 -247 373 -246
rect 373 -247 374 -246
rect 374 -247 375 -246
rect 375 -247 376 -246
rect 376 -247 377 -246
rect 377 -247 378 -246
rect 378 -247 379 -246
rect 379 -247 380 -246
rect 380 -247 381 -246
rect 381 -247 382 -246
rect 382 -247 383 -246
rect 383 -247 384 -246
rect 384 -247 385 -246
rect 385 -247 386 -246
rect 386 -247 387 -246
rect 387 -247 388 -246
rect 388 -247 389 -246
rect 389 -247 390 -246
rect 390 -247 391 -246
rect 391 -247 392 -246
rect 392 -247 393 -246
rect 393 -247 394 -246
rect 394 -247 395 -246
rect 395 -247 396 -246
rect 396 -247 397 -246
rect 397 -247 398 -246
rect 398 -247 399 -246
rect 399 -247 400 -246
rect 400 -247 401 -246
rect 401 -247 402 -246
rect 402 -247 403 -246
rect 403 -247 404 -246
rect 404 -247 405 -246
rect 405 -247 406 -246
rect 406 -247 407 -246
rect 407 -247 408 -246
rect 408 -247 409 -246
rect 409 -247 410 -246
rect 410 -247 411 -246
rect 411 -247 412 -246
rect 412 -247 413 -246
rect 413 -247 414 -246
rect 414 -247 415 -246
rect 415 -247 416 -246
rect 416 -247 417 -246
rect 417 -247 418 -246
rect 418 -247 419 -246
rect 419 -247 420 -246
rect 420 -247 421 -246
rect 421 -247 422 -246
rect 422 -247 423 -246
rect 423 -247 424 -246
rect 424 -247 425 -246
rect 425 -247 426 -246
rect 426 -247 427 -246
rect 427 -247 428 -246
rect 428 -247 429 -246
rect 429 -247 430 -246
rect 430 -247 431 -246
rect 431 -247 432 -246
rect 432 -247 433 -246
rect 433 -247 434 -246
rect 434 -247 435 -246
rect 435 -247 436 -246
rect 436 -247 437 -246
rect 437 -247 438 -246
rect 438 -247 439 -246
rect 439 -247 440 -246
rect 440 -247 441 -246
rect 441 -247 442 -246
rect 442 -247 443 -246
rect 443 -247 444 -246
rect 444 -247 445 -246
rect 445 -247 446 -246
rect 446 -247 447 -246
rect 447 -247 448 -246
rect 448 -247 449 -246
rect 449 -247 450 -246
rect 450 -247 451 -246
rect 451 -247 452 -246
rect 452 -247 453 -246
rect 453 -247 454 -246
rect 454 -247 455 -246
rect 455 -247 456 -246
rect 456 -247 457 -246
rect 457 -247 458 -246
rect 458 -247 459 -246
rect 459 -247 460 -246
rect 460 -247 461 -246
rect 461 -247 462 -246
rect 462 -247 463 -246
rect 463 -247 464 -246
rect 464 -247 465 -246
rect 465 -247 466 -246
rect 466 -247 467 -246
rect 467 -247 468 -246
rect 468 -247 469 -246
rect 469 -247 470 -246
rect 470 -247 471 -246
rect 471 -247 472 -246
rect 472 -247 473 -246
rect 473 -247 474 -246
rect 474 -247 475 -246
rect 475 -247 476 -246
rect 476 -247 477 -246
rect 477 -247 478 -246
rect 478 -247 479 -246
rect 479 -247 480 -246
rect 2 -248 3 -247
rect 3 -248 4 -247
rect 4 -248 5 -247
rect 5 -248 6 -247
rect 6 -248 7 -247
rect 7 -248 8 -247
rect 8 -248 9 -247
rect 9 -248 10 -247
rect 10 -248 11 -247
rect 11 -248 12 -247
rect 12 -248 13 -247
rect 13 -248 14 -247
rect 14 -248 15 -247
rect 15 -248 16 -247
rect 16 -248 17 -247
rect 17 -248 18 -247
rect 18 -248 19 -247
rect 19 -248 20 -247
rect 20 -248 21 -247
rect 21 -248 22 -247
rect 22 -248 23 -247
rect 23 -248 24 -247
rect 24 -248 25 -247
rect 25 -248 26 -247
rect 26 -248 27 -247
rect 27 -248 28 -247
rect 28 -248 29 -247
rect 29 -248 30 -247
rect 30 -248 31 -247
rect 31 -248 32 -247
rect 32 -248 33 -247
rect 33 -248 34 -247
rect 34 -248 35 -247
rect 35 -248 36 -247
rect 36 -248 37 -247
rect 37 -248 38 -247
rect 38 -248 39 -247
rect 39 -248 40 -247
rect 40 -248 41 -247
rect 41 -248 42 -247
rect 42 -248 43 -247
rect 43 -248 44 -247
rect 44 -248 45 -247
rect 45 -248 46 -247
rect 46 -248 47 -247
rect 47 -248 48 -247
rect 48 -248 49 -247
rect 49 -248 50 -247
rect 50 -248 51 -247
rect 51 -248 52 -247
rect 52 -248 53 -247
rect 53 -248 54 -247
rect 54 -248 55 -247
rect 55 -248 56 -247
rect 56 -248 57 -247
rect 57 -248 58 -247
rect 58 -248 59 -247
rect 59 -248 60 -247
rect 60 -248 61 -247
rect 61 -248 62 -247
rect 62 -248 63 -247
rect 63 -248 64 -247
rect 64 -248 65 -247
rect 65 -248 66 -247
rect 66 -248 67 -247
rect 67 -248 68 -247
rect 68 -248 69 -247
rect 69 -248 70 -247
rect 70 -248 71 -247
rect 71 -248 72 -247
rect 72 -248 73 -247
rect 73 -248 74 -247
rect 74 -248 75 -247
rect 75 -248 76 -247
rect 76 -248 77 -247
rect 77 -248 78 -247
rect 78 -248 79 -247
rect 79 -248 80 -247
rect 80 -248 81 -247
rect 81 -248 82 -247
rect 82 -248 83 -247
rect 83 -248 84 -247
rect 84 -248 85 -247
rect 85 -248 86 -247
rect 86 -248 87 -247
rect 87 -248 88 -247
rect 88 -248 89 -247
rect 89 -248 90 -247
rect 90 -248 91 -247
rect 91 -248 92 -247
rect 92 -248 93 -247
rect 93 -248 94 -247
rect 94 -248 95 -247
rect 95 -248 96 -247
rect 96 -248 97 -247
rect 97 -248 98 -247
rect 98 -248 99 -247
rect 99 -248 100 -247
rect 100 -248 101 -247
rect 101 -248 102 -247
rect 102 -248 103 -247
rect 103 -248 104 -247
rect 104 -248 105 -247
rect 105 -248 106 -247
rect 106 -248 107 -247
rect 107 -248 108 -247
rect 108 -248 109 -247
rect 109 -248 110 -247
rect 110 -248 111 -247
rect 111 -248 112 -247
rect 112 -248 113 -247
rect 113 -248 114 -247
rect 114 -248 115 -247
rect 115 -248 116 -247
rect 116 -248 117 -247
rect 117 -248 118 -247
rect 118 -248 119 -247
rect 119 -248 120 -247
rect 120 -248 121 -247
rect 121 -248 122 -247
rect 122 -248 123 -247
rect 123 -248 124 -247
rect 124 -248 125 -247
rect 125 -248 126 -247
rect 126 -248 127 -247
rect 127 -248 128 -247
rect 128 -248 129 -247
rect 129 -248 130 -247
rect 130 -248 131 -247
rect 131 -248 132 -247
rect 132 -248 133 -247
rect 133 -248 134 -247
rect 134 -248 135 -247
rect 135 -248 136 -247
rect 136 -248 137 -247
rect 137 -248 138 -247
rect 138 -248 139 -247
rect 139 -248 140 -247
rect 140 -248 141 -247
rect 141 -248 142 -247
rect 142 -248 143 -247
rect 143 -248 144 -247
rect 144 -248 145 -247
rect 145 -248 146 -247
rect 146 -248 147 -247
rect 147 -248 148 -247
rect 148 -248 149 -247
rect 149 -248 150 -247
rect 150 -248 151 -247
rect 151 -248 152 -247
rect 152 -248 153 -247
rect 153 -248 154 -247
rect 154 -248 155 -247
rect 155 -248 156 -247
rect 156 -248 157 -247
rect 157 -248 158 -247
rect 158 -248 159 -247
rect 159 -248 160 -247
rect 160 -248 161 -247
rect 161 -248 162 -247
rect 162 -248 163 -247
rect 163 -248 164 -247
rect 164 -248 165 -247
rect 165 -248 166 -247
rect 166 -248 167 -247
rect 167 -248 168 -247
rect 168 -248 169 -247
rect 169 -248 170 -247
rect 170 -248 171 -247
rect 171 -248 172 -247
rect 172 -248 173 -247
rect 173 -248 174 -247
rect 174 -248 175 -247
rect 175 -248 176 -247
rect 176 -248 177 -247
rect 177 -248 178 -247
rect 178 -248 179 -247
rect 179 -248 180 -247
rect 180 -248 181 -247
rect 181 -248 182 -247
rect 182 -248 183 -247
rect 183 -248 184 -247
rect 184 -248 185 -247
rect 185 -248 186 -247
rect 186 -248 187 -247
rect 187 -248 188 -247
rect 188 -248 189 -247
rect 189 -248 190 -247
rect 190 -248 191 -247
rect 191 -248 192 -247
rect 192 -248 193 -247
rect 193 -248 194 -247
rect 194 -248 195 -247
rect 195 -248 196 -247
rect 196 -248 197 -247
rect 197 -248 198 -247
rect 198 -248 199 -247
rect 199 -248 200 -247
rect 200 -248 201 -247
rect 201 -248 202 -247
rect 202 -248 203 -247
rect 203 -248 204 -247
rect 204 -248 205 -247
rect 205 -248 206 -247
rect 206 -248 207 -247
rect 207 -248 208 -247
rect 208 -248 209 -247
rect 209 -248 210 -247
rect 210 -248 211 -247
rect 211 -248 212 -247
rect 212 -248 213 -247
rect 213 -248 214 -247
rect 214 -248 215 -247
rect 215 -248 216 -247
rect 216 -248 217 -247
rect 217 -248 218 -247
rect 218 -248 219 -247
rect 219 -248 220 -247
rect 220 -248 221 -247
rect 221 -248 222 -247
rect 222 -248 223 -247
rect 223 -248 224 -247
rect 224 -248 225 -247
rect 225 -248 226 -247
rect 226 -248 227 -247
rect 227 -248 228 -247
rect 228 -248 229 -247
rect 229 -248 230 -247
rect 230 -248 231 -247
rect 231 -248 232 -247
rect 232 -248 233 -247
rect 233 -248 234 -247
rect 234 -248 235 -247
rect 235 -248 236 -247
rect 236 -248 237 -247
rect 237 -248 238 -247
rect 238 -248 239 -247
rect 239 -248 240 -247
rect 240 -248 241 -247
rect 241 -248 242 -247
rect 242 -248 243 -247
rect 243 -248 244 -247
rect 244 -248 245 -247
rect 245 -248 246 -247
rect 246 -248 247 -247
rect 247 -248 248 -247
rect 248 -248 249 -247
rect 249 -248 250 -247
rect 250 -248 251 -247
rect 251 -248 252 -247
rect 252 -248 253 -247
rect 253 -248 254 -247
rect 254 -248 255 -247
rect 255 -248 256 -247
rect 256 -248 257 -247
rect 257 -248 258 -247
rect 258 -248 259 -247
rect 259 -248 260 -247
rect 260 -248 261 -247
rect 261 -248 262 -247
rect 262 -248 263 -247
rect 263 -248 264 -247
rect 264 -248 265 -247
rect 265 -248 266 -247
rect 266 -248 267 -247
rect 267 -248 268 -247
rect 268 -248 269 -247
rect 269 -248 270 -247
rect 270 -248 271 -247
rect 271 -248 272 -247
rect 272 -248 273 -247
rect 273 -248 274 -247
rect 274 -248 275 -247
rect 275 -248 276 -247
rect 276 -248 277 -247
rect 277 -248 278 -247
rect 278 -248 279 -247
rect 279 -248 280 -247
rect 280 -248 281 -247
rect 281 -248 282 -247
rect 282 -248 283 -247
rect 283 -248 284 -247
rect 284 -248 285 -247
rect 285 -248 286 -247
rect 286 -248 287 -247
rect 287 -248 288 -247
rect 288 -248 289 -247
rect 289 -248 290 -247
rect 290 -248 291 -247
rect 291 -248 292 -247
rect 292 -248 293 -247
rect 293 -248 294 -247
rect 294 -248 295 -247
rect 295 -248 296 -247
rect 296 -248 297 -247
rect 297 -248 298 -247
rect 298 -248 299 -247
rect 299 -248 300 -247
rect 300 -248 301 -247
rect 301 -248 302 -247
rect 302 -248 303 -247
rect 303 -248 304 -247
rect 304 -248 305 -247
rect 305 -248 306 -247
rect 306 -248 307 -247
rect 307 -248 308 -247
rect 308 -248 309 -247
rect 309 -248 310 -247
rect 310 -248 311 -247
rect 311 -248 312 -247
rect 312 -248 313 -247
rect 313 -248 314 -247
rect 314 -248 315 -247
rect 315 -248 316 -247
rect 316 -248 317 -247
rect 317 -248 318 -247
rect 318 -248 319 -247
rect 319 -248 320 -247
rect 320 -248 321 -247
rect 321 -248 322 -247
rect 322 -248 323 -247
rect 323 -248 324 -247
rect 324 -248 325 -247
rect 325 -248 326 -247
rect 326 -248 327 -247
rect 327 -248 328 -247
rect 328 -248 329 -247
rect 329 -248 330 -247
rect 330 -248 331 -247
rect 331 -248 332 -247
rect 332 -248 333 -247
rect 333 -248 334 -247
rect 334 -248 335 -247
rect 335 -248 336 -247
rect 336 -248 337 -247
rect 337 -248 338 -247
rect 338 -248 339 -247
rect 339 -248 340 -247
rect 340 -248 341 -247
rect 341 -248 342 -247
rect 342 -248 343 -247
rect 343 -248 344 -247
rect 344 -248 345 -247
rect 345 -248 346 -247
rect 346 -248 347 -247
rect 347 -248 348 -247
rect 348 -248 349 -247
rect 349 -248 350 -247
rect 350 -248 351 -247
rect 351 -248 352 -247
rect 352 -248 353 -247
rect 353 -248 354 -247
rect 354 -248 355 -247
rect 355 -248 356 -247
rect 356 -248 357 -247
rect 357 -248 358 -247
rect 358 -248 359 -247
rect 359 -248 360 -247
rect 360 -248 361 -247
rect 361 -248 362 -247
rect 362 -248 363 -247
rect 363 -248 364 -247
rect 364 -248 365 -247
rect 365 -248 366 -247
rect 366 -248 367 -247
rect 367 -248 368 -247
rect 368 -248 369 -247
rect 369 -248 370 -247
rect 370 -248 371 -247
rect 371 -248 372 -247
rect 372 -248 373 -247
rect 373 -248 374 -247
rect 374 -248 375 -247
rect 375 -248 376 -247
rect 376 -248 377 -247
rect 377 -248 378 -247
rect 378 -248 379 -247
rect 379 -248 380 -247
rect 380 -248 381 -247
rect 381 -248 382 -247
rect 382 -248 383 -247
rect 383 -248 384 -247
rect 384 -248 385 -247
rect 385 -248 386 -247
rect 386 -248 387 -247
rect 387 -248 388 -247
rect 388 -248 389 -247
rect 389 -248 390 -247
rect 390 -248 391 -247
rect 391 -248 392 -247
rect 392 -248 393 -247
rect 393 -248 394 -247
rect 394 -248 395 -247
rect 395 -248 396 -247
rect 396 -248 397 -247
rect 397 -248 398 -247
rect 398 -248 399 -247
rect 399 -248 400 -247
rect 400 -248 401 -247
rect 401 -248 402 -247
rect 402 -248 403 -247
rect 403 -248 404 -247
rect 404 -248 405 -247
rect 405 -248 406 -247
rect 406 -248 407 -247
rect 407 -248 408 -247
rect 408 -248 409 -247
rect 409 -248 410 -247
rect 410 -248 411 -247
rect 411 -248 412 -247
rect 412 -248 413 -247
rect 413 -248 414 -247
rect 414 -248 415 -247
rect 415 -248 416 -247
rect 416 -248 417 -247
rect 417 -248 418 -247
rect 418 -248 419 -247
rect 419 -248 420 -247
rect 420 -248 421 -247
rect 421 -248 422 -247
rect 422 -248 423 -247
rect 423 -248 424 -247
rect 424 -248 425 -247
rect 425 -248 426 -247
rect 426 -248 427 -247
rect 427 -248 428 -247
rect 428 -248 429 -247
rect 429 -248 430 -247
rect 430 -248 431 -247
rect 431 -248 432 -247
rect 432 -248 433 -247
rect 433 -248 434 -247
rect 434 -248 435 -247
rect 435 -248 436 -247
rect 436 -248 437 -247
rect 437 -248 438 -247
rect 438 -248 439 -247
rect 439 -248 440 -247
rect 440 -248 441 -247
rect 441 -248 442 -247
rect 442 -248 443 -247
rect 443 -248 444 -247
rect 444 -248 445 -247
rect 445 -248 446 -247
rect 446 -248 447 -247
rect 447 -248 448 -247
rect 448 -248 449 -247
rect 449 -248 450 -247
rect 450 -248 451 -247
rect 451 -248 452 -247
rect 452 -248 453 -247
rect 453 -248 454 -247
rect 454 -248 455 -247
rect 455 -248 456 -247
rect 456 -248 457 -247
rect 457 -248 458 -247
rect 458 -248 459 -247
rect 459 -248 460 -247
rect 460 -248 461 -247
rect 461 -248 462 -247
rect 462 -248 463 -247
rect 463 -248 464 -247
rect 464 -248 465 -247
rect 465 -248 466 -247
rect 466 -248 467 -247
rect 467 -248 468 -247
rect 468 -248 469 -247
rect 469 -248 470 -247
rect 470 -248 471 -247
rect 471 -248 472 -247
rect 472 -248 473 -247
rect 473 -248 474 -247
rect 474 -248 475 -247
rect 475 -248 476 -247
rect 476 -248 477 -247
rect 477 -248 478 -247
rect 478 -248 479 -247
rect 479 -248 480 -247
rect 2 -249 3 -248
rect 3 -249 4 -248
rect 4 -249 5 -248
rect 5 -249 6 -248
rect 6 -249 7 -248
rect 7 -249 8 -248
rect 8 -249 9 -248
rect 9 -249 10 -248
rect 10 -249 11 -248
rect 11 -249 12 -248
rect 12 -249 13 -248
rect 13 -249 14 -248
rect 14 -249 15 -248
rect 15 -249 16 -248
rect 16 -249 17 -248
rect 17 -249 18 -248
rect 18 -249 19 -248
rect 19 -249 20 -248
rect 20 -249 21 -248
rect 21 -249 22 -248
rect 22 -249 23 -248
rect 23 -249 24 -248
rect 24 -249 25 -248
rect 25 -249 26 -248
rect 26 -249 27 -248
rect 27 -249 28 -248
rect 28 -249 29 -248
rect 29 -249 30 -248
rect 30 -249 31 -248
rect 31 -249 32 -248
rect 32 -249 33 -248
rect 33 -249 34 -248
rect 34 -249 35 -248
rect 35 -249 36 -248
rect 36 -249 37 -248
rect 37 -249 38 -248
rect 38 -249 39 -248
rect 39 -249 40 -248
rect 40 -249 41 -248
rect 41 -249 42 -248
rect 42 -249 43 -248
rect 43 -249 44 -248
rect 44 -249 45 -248
rect 45 -249 46 -248
rect 46 -249 47 -248
rect 47 -249 48 -248
rect 48 -249 49 -248
rect 49 -249 50 -248
rect 50 -249 51 -248
rect 51 -249 52 -248
rect 52 -249 53 -248
rect 53 -249 54 -248
rect 54 -249 55 -248
rect 55 -249 56 -248
rect 56 -249 57 -248
rect 57 -249 58 -248
rect 58 -249 59 -248
rect 59 -249 60 -248
rect 60 -249 61 -248
rect 61 -249 62 -248
rect 62 -249 63 -248
rect 63 -249 64 -248
rect 64 -249 65 -248
rect 65 -249 66 -248
rect 66 -249 67 -248
rect 67 -249 68 -248
rect 68 -249 69 -248
rect 69 -249 70 -248
rect 70 -249 71 -248
rect 71 -249 72 -248
rect 72 -249 73 -248
rect 73 -249 74 -248
rect 74 -249 75 -248
rect 75 -249 76 -248
rect 76 -249 77 -248
rect 77 -249 78 -248
rect 78 -249 79 -248
rect 79 -249 80 -248
rect 80 -249 81 -248
rect 81 -249 82 -248
rect 82 -249 83 -248
rect 83 -249 84 -248
rect 84 -249 85 -248
rect 85 -249 86 -248
rect 86 -249 87 -248
rect 87 -249 88 -248
rect 88 -249 89 -248
rect 89 -249 90 -248
rect 90 -249 91 -248
rect 91 -249 92 -248
rect 92 -249 93 -248
rect 93 -249 94 -248
rect 94 -249 95 -248
rect 95 -249 96 -248
rect 96 -249 97 -248
rect 97 -249 98 -248
rect 98 -249 99 -248
rect 99 -249 100 -248
rect 100 -249 101 -248
rect 101 -249 102 -248
rect 102 -249 103 -248
rect 103 -249 104 -248
rect 104 -249 105 -248
rect 105 -249 106 -248
rect 106 -249 107 -248
rect 107 -249 108 -248
rect 108 -249 109 -248
rect 109 -249 110 -248
rect 110 -249 111 -248
rect 111 -249 112 -248
rect 112 -249 113 -248
rect 113 -249 114 -248
rect 114 -249 115 -248
rect 115 -249 116 -248
rect 116 -249 117 -248
rect 117 -249 118 -248
rect 118 -249 119 -248
rect 119 -249 120 -248
rect 120 -249 121 -248
rect 121 -249 122 -248
rect 122 -249 123 -248
rect 123 -249 124 -248
rect 124 -249 125 -248
rect 125 -249 126 -248
rect 126 -249 127 -248
rect 127 -249 128 -248
rect 128 -249 129 -248
rect 129 -249 130 -248
rect 130 -249 131 -248
rect 131 -249 132 -248
rect 132 -249 133 -248
rect 133 -249 134 -248
rect 134 -249 135 -248
rect 135 -249 136 -248
rect 136 -249 137 -248
rect 137 -249 138 -248
rect 138 -249 139 -248
rect 139 -249 140 -248
rect 140 -249 141 -248
rect 141 -249 142 -248
rect 142 -249 143 -248
rect 143 -249 144 -248
rect 144 -249 145 -248
rect 145 -249 146 -248
rect 146 -249 147 -248
rect 147 -249 148 -248
rect 148 -249 149 -248
rect 149 -249 150 -248
rect 150 -249 151 -248
rect 151 -249 152 -248
rect 152 -249 153 -248
rect 153 -249 154 -248
rect 154 -249 155 -248
rect 155 -249 156 -248
rect 156 -249 157 -248
rect 157 -249 158 -248
rect 158 -249 159 -248
rect 159 -249 160 -248
rect 160 -249 161 -248
rect 161 -249 162 -248
rect 162 -249 163 -248
rect 163 -249 164 -248
rect 164 -249 165 -248
rect 165 -249 166 -248
rect 166 -249 167 -248
rect 167 -249 168 -248
rect 168 -249 169 -248
rect 169 -249 170 -248
rect 170 -249 171 -248
rect 171 -249 172 -248
rect 172 -249 173 -248
rect 173 -249 174 -248
rect 174 -249 175 -248
rect 175 -249 176 -248
rect 176 -249 177 -248
rect 177 -249 178 -248
rect 178 -249 179 -248
rect 179 -249 180 -248
rect 180 -249 181 -248
rect 181 -249 182 -248
rect 182 -249 183 -248
rect 183 -249 184 -248
rect 184 -249 185 -248
rect 185 -249 186 -248
rect 186 -249 187 -248
rect 187 -249 188 -248
rect 188 -249 189 -248
rect 189 -249 190 -248
rect 190 -249 191 -248
rect 191 -249 192 -248
rect 192 -249 193 -248
rect 193 -249 194 -248
rect 194 -249 195 -248
rect 195 -249 196 -248
rect 196 -249 197 -248
rect 197 -249 198 -248
rect 198 -249 199 -248
rect 199 -249 200 -248
rect 200 -249 201 -248
rect 201 -249 202 -248
rect 202 -249 203 -248
rect 203 -249 204 -248
rect 204 -249 205 -248
rect 205 -249 206 -248
rect 206 -249 207 -248
rect 207 -249 208 -248
rect 208 -249 209 -248
rect 209 -249 210 -248
rect 210 -249 211 -248
rect 211 -249 212 -248
rect 212 -249 213 -248
rect 213 -249 214 -248
rect 214 -249 215 -248
rect 215 -249 216 -248
rect 216 -249 217 -248
rect 217 -249 218 -248
rect 218 -249 219 -248
rect 219 -249 220 -248
rect 220 -249 221 -248
rect 221 -249 222 -248
rect 222 -249 223 -248
rect 223 -249 224 -248
rect 224 -249 225 -248
rect 225 -249 226 -248
rect 226 -249 227 -248
rect 227 -249 228 -248
rect 228 -249 229 -248
rect 229 -249 230 -248
rect 230 -249 231 -248
rect 231 -249 232 -248
rect 232 -249 233 -248
rect 233 -249 234 -248
rect 234 -249 235 -248
rect 235 -249 236 -248
rect 236 -249 237 -248
rect 237 -249 238 -248
rect 238 -249 239 -248
rect 239 -249 240 -248
rect 240 -249 241 -248
rect 241 -249 242 -248
rect 242 -249 243 -248
rect 243 -249 244 -248
rect 244 -249 245 -248
rect 245 -249 246 -248
rect 246 -249 247 -248
rect 247 -249 248 -248
rect 248 -249 249 -248
rect 249 -249 250 -248
rect 250 -249 251 -248
rect 251 -249 252 -248
rect 252 -249 253 -248
rect 253 -249 254 -248
rect 254 -249 255 -248
rect 255 -249 256 -248
rect 256 -249 257 -248
rect 257 -249 258 -248
rect 258 -249 259 -248
rect 259 -249 260 -248
rect 260 -249 261 -248
rect 261 -249 262 -248
rect 262 -249 263 -248
rect 263 -249 264 -248
rect 264 -249 265 -248
rect 265 -249 266 -248
rect 266 -249 267 -248
rect 267 -249 268 -248
rect 268 -249 269 -248
rect 269 -249 270 -248
rect 270 -249 271 -248
rect 271 -249 272 -248
rect 272 -249 273 -248
rect 273 -249 274 -248
rect 274 -249 275 -248
rect 275 -249 276 -248
rect 276 -249 277 -248
rect 277 -249 278 -248
rect 278 -249 279 -248
rect 279 -249 280 -248
rect 280 -249 281 -248
rect 281 -249 282 -248
rect 282 -249 283 -248
rect 283 -249 284 -248
rect 284 -249 285 -248
rect 285 -249 286 -248
rect 286 -249 287 -248
rect 287 -249 288 -248
rect 288 -249 289 -248
rect 289 -249 290 -248
rect 290 -249 291 -248
rect 291 -249 292 -248
rect 292 -249 293 -248
rect 293 -249 294 -248
rect 294 -249 295 -248
rect 295 -249 296 -248
rect 296 -249 297 -248
rect 297 -249 298 -248
rect 298 -249 299 -248
rect 299 -249 300 -248
rect 300 -249 301 -248
rect 301 -249 302 -248
rect 302 -249 303 -248
rect 303 -249 304 -248
rect 304 -249 305 -248
rect 305 -249 306 -248
rect 306 -249 307 -248
rect 307 -249 308 -248
rect 308 -249 309 -248
rect 309 -249 310 -248
rect 310 -249 311 -248
rect 311 -249 312 -248
rect 312 -249 313 -248
rect 313 -249 314 -248
rect 314 -249 315 -248
rect 315 -249 316 -248
rect 316 -249 317 -248
rect 317 -249 318 -248
rect 318 -249 319 -248
rect 319 -249 320 -248
rect 320 -249 321 -248
rect 321 -249 322 -248
rect 322 -249 323 -248
rect 323 -249 324 -248
rect 324 -249 325 -248
rect 325 -249 326 -248
rect 326 -249 327 -248
rect 327 -249 328 -248
rect 328 -249 329 -248
rect 329 -249 330 -248
rect 330 -249 331 -248
rect 331 -249 332 -248
rect 332 -249 333 -248
rect 333 -249 334 -248
rect 334 -249 335 -248
rect 335 -249 336 -248
rect 336 -249 337 -248
rect 337 -249 338 -248
rect 338 -249 339 -248
rect 339 -249 340 -248
rect 340 -249 341 -248
rect 341 -249 342 -248
rect 342 -249 343 -248
rect 343 -249 344 -248
rect 344 -249 345 -248
rect 345 -249 346 -248
rect 346 -249 347 -248
rect 347 -249 348 -248
rect 348 -249 349 -248
rect 349 -249 350 -248
rect 350 -249 351 -248
rect 351 -249 352 -248
rect 352 -249 353 -248
rect 353 -249 354 -248
rect 354 -249 355 -248
rect 355 -249 356 -248
rect 356 -249 357 -248
rect 357 -249 358 -248
rect 358 -249 359 -248
rect 359 -249 360 -248
rect 360 -249 361 -248
rect 361 -249 362 -248
rect 362 -249 363 -248
rect 363 -249 364 -248
rect 364 -249 365 -248
rect 365 -249 366 -248
rect 366 -249 367 -248
rect 367 -249 368 -248
rect 368 -249 369 -248
rect 369 -249 370 -248
rect 370 -249 371 -248
rect 371 -249 372 -248
rect 372 -249 373 -248
rect 373 -249 374 -248
rect 374 -249 375 -248
rect 375 -249 376 -248
rect 376 -249 377 -248
rect 377 -249 378 -248
rect 378 -249 379 -248
rect 379 -249 380 -248
rect 380 -249 381 -248
rect 381 -249 382 -248
rect 382 -249 383 -248
rect 383 -249 384 -248
rect 384 -249 385 -248
rect 385 -249 386 -248
rect 386 -249 387 -248
rect 387 -249 388 -248
rect 388 -249 389 -248
rect 389 -249 390 -248
rect 390 -249 391 -248
rect 391 -249 392 -248
rect 392 -249 393 -248
rect 393 -249 394 -248
rect 394 -249 395 -248
rect 395 -249 396 -248
rect 396 -249 397 -248
rect 397 -249 398 -248
rect 398 -249 399 -248
rect 399 -249 400 -248
rect 400 -249 401 -248
rect 401 -249 402 -248
rect 402 -249 403 -248
rect 403 -249 404 -248
rect 404 -249 405 -248
rect 405 -249 406 -248
rect 406 -249 407 -248
rect 407 -249 408 -248
rect 408 -249 409 -248
rect 409 -249 410 -248
rect 410 -249 411 -248
rect 411 -249 412 -248
rect 412 -249 413 -248
rect 413 -249 414 -248
rect 414 -249 415 -248
rect 415 -249 416 -248
rect 416 -249 417 -248
rect 417 -249 418 -248
rect 418 -249 419 -248
rect 419 -249 420 -248
rect 420 -249 421 -248
rect 421 -249 422 -248
rect 422 -249 423 -248
rect 423 -249 424 -248
rect 424 -249 425 -248
rect 425 -249 426 -248
rect 426 -249 427 -248
rect 427 -249 428 -248
rect 428 -249 429 -248
rect 429 -249 430 -248
rect 430 -249 431 -248
rect 431 -249 432 -248
rect 432 -249 433 -248
rect 433 -249 434 -248
rect 434 -249 435 -248
rect 435 -249 436 -248
rect 436 -249 437 -248
rect 437 -249 438 -248
rect 438 -249 439 -248
rect 439 -249 440 -248
rect 440 -249 441 -248
rect 441 -249 442 -248
rect 442 -249 443 -248
rect 443 -249 444 -248
rect 444 -249 445 -248
rect 445 -249 446 -248
rect 446 -249 447 -248
rect 447 -249 448 -248
rect 448 -249 449 -248
rect 449 -249 450 -248
rect 450 -249 451 -248
rect 451 -249 452 -248
rect 452 -249 453 -248
rect 453 -249 454 -248
rect 454 -249 455 -248
rect 455 -249 456 -248
rect 456 -249 457 -248
rect 457 -249 458 -248
rect 458 -249 459 -248
rect 459 -249 460 -248
rect 460 -249 461 -248
rect 461 -249 462 -248
rect 462 -249 463 -248
rect 463 -249 464 -248
rect 464 -249 465 -248
rect 465 -249 466 -248
rect 466 -249 467 -248
rect 467 -249 468 -248
rect 468 -249 469 -248
rect 469 -249 470 -248
rect 470 -249 471 -248
rect 471 -249 472 -248
rect 472 -249 473 -248
rect 473 -249 474 -248
rect 474 -249 475 -248
rect 475 -249 476 -248
rect 476 -249 477 -248
rect 477 -249 478 -248
rect 478 -249 479 -248
rect 479 -249 480 -248
rect 2 -250 3 -249
rect 3 -250 4 -249
rect 4 -250 5 -249
rect 5 -250 6 -249
rect 6 -250 7 -249
rect 7 -250 8 -249
rect 8 -250 9 -249
rect 9 -250 10 -249
rect 10 -250 11 -249
rect 11 -250 12 -249
rect 12 -250 13 -249
rect 13 -250 14 -249
rect 14 -250 15 -249
rect 15 -250 16 -249
rect 16 -250 17 -249
rect 17 -250 18 -249
rect 18 -250 19 -249
rect 19 -250 20 -249
rect 20 -250 21 -249
rect 21 -250 22 -249
rect 22 -250 23 -249
rect 23 -250 24 -249
rect 24 -250 25 -249
rect 25 -250 26 -249
rect 26 -250 27 -249
rect 27 -250 28 -249
rect 28 -250 29 -249
rect 29 -250 30 -249
rect 30 -250 31 -249
rect 31 -250 32 -249
rect 32 -250 33 -249
rect 33 -250 34 -249
rect 34 -250 35 -249
rect 35 -250 36 -249
rect 36 -250 37 -249
rect 37 -250 38 -249
rect 38 -250 39 -249
rect 39 -250 40 -249
rect 40 -250 41 -249
rect 41 -250 42 -249
rect 42 -250 43 -249
rect 43 -250 44 -249
rect 44 -250 45 -249
rect 45 -250 46 -249
rect 46 -250 47 -249
rect 47 -250 48 -249
rect 48 -250 49 -249
rect 49 -250 50 -249
rect 50 -250 51 -249
rect 51 -250 52 -249
rect 52 -250 53 -249
rect 53 -250 54 -249
rect 54 -250 55 -249
rect 55 -250 56 -249
rect 56 -250 57 -249
rect 57 -250 58 -249
rect 58 -250 59 -249
rect 59 -250 60 -249
rect 60 -250 61 -249
rect 61 -250 62 -249
rect 62 -250 63 -249
rect 63 -250 64 -249
rect 64 -250 65 -249
rect 65 -250 66 -249
rect 66 -250 67 -249
rect 67 -250 68 -249
rect 68 -250 69 -249
rect 69 -250 70 -249
rect 70 -250 71 -249
rect 71 -250 72 -249
rect 72 -250 73 -249
rect 73 -250 74 -249
rect 74 -250 75 -249
rect 75 -250 76 -249
rect 76 -250 77 -249
rect 77 -250 78 -249
rect 78 -250 79 -249
rect 79 -250 80 -249
rect 80 -250 81 -249
rect 81 -250 82 -249
rect 82 -250 83 -249
rect 83 -250 84 -249
rect 84 -250 85 -249
rect 85 -250 86 -249
rect 86 -250 87 -249
rect 87 -250 88 -249
rect 88 -250 89 -249
rect 89 -250 90 -249
rect 90 -250 91 -249
rect 91 -250 92 -249
rect 92 -250 93 -249
rect 93 -250 94 -249
rect 94 -250 95 -249
rect 95 -250 96 -249
rect 96 -250 97 -249
rect 97 -250 98 -249
rect 98 -250 99 -249
rect 99 -250 100 -249
rect 100 -250 101 -249
rect 101 -250 102 -249
rect 102 -250 103 -249
rect 103 -250 104 -249
rect 104 -250 105 -249
rect 105 -250 106 -249
rect 106 -250 107 -249
rect 107 -250 108 -249
rect 108 -250 109 -249
rect 109 -250 110 -249
rect 110 -250 111 -249
rect 111 -250 112 -249
rect 112 -250 113 -249
rect 113 -250 114 -249
rect 114 -250 115 -249
rect 115 -250 116 -249
rect 116 -250 117 -249
rect 117 -250 118 -249
rect 118 -250 119 -249
rect 119 -250 120 -249
rect 120 -250 121 -249
rect 121 -250 122 -249
rect 122 -250 123 -249
rect 123 -250 124 -249
rect 124 -250 125 -249
rect 125 -250 126 -249
rect 126 -250 127 -249
rect 127 -250 128 -249
rect 128 -250 129 -249
rect 129 -250 130 -249
rect 130 -250 131 -249
rect 131 -250 132 -249
rect 132 -250 133 -249
rect 133 -250 134 -249
rect 134 -250 135 -249
rect 135 -250 136 -249
rect 136 -250 137 -249
rect 137 -250 138 -249
rect 138 -250 139 -249
rect 139 -250 140 -249
rect 140 -250 141 -249
rect 141 -250 142 -249
rect 142 -250 143 -249
rect 143 -250 144 -249
rect 144 -250 145 -249
rect 145 -250 146 -249
rect 146 -250 147 -249
rect 147 -250 148 -249
rect 148 -250 149 -249
rect 149 -250 150 -249
rect 150 -250 151 -249
rect 151 -250 152 -249
rect 152 -250 153 -249
rect 153 -250 154 -249
rect 154 -250 155 -249
rect 155 -250 156 -249
rect 156 -250 157 -249
rect 157 -250 158 -249
rect 158 -250 159 -249
rect 159 -250 160 -249
rect 160 -250 161 -249
rect 161 -250 162 -249
rect 162 -250 163 -249
rect 163 -250 164 -249
rect 164 -250 165 -249
rect 165 -250 166 -249
rect 166 -250 167 -249
rect 167 -250 168 -249
rect 168 -250 169 -249
rect 169 -250 170 -249
rect 170 -250 171 -249
rect 171 -250 172 -249
rect 172 -250 173 -249
rect 173 -250 174 -249
rect 174 -250 175 -249
rect 175 -250 176 -249
rect 176 -250 177 -249
rect 177 -250 178 -249
rect 178 -250 179 -249
rect 179 -250 180 -249
rect 180 -250 181 -249
rect 181 -250 182 -249
rect 182 -250 183 -249
rect 183 -250 184 -249
rect 184 -250 185 -249
rect 185 -250 186 -249
rect 186 -250 187 -249
rect 187 -250 188 -249
rect 188 -250 189 -249
rect 189 -250 190 -249
rect 190 -250 191 -249
rect 191 -250 192 -249
rect 192 -250 193 -249
rect 193 -250 194 -249
rect 194 -250 195 -249
rect 195 -250 196 -249
rect 196 -250 197 -249
rect 197 -250 198 -249
rect 198 -250 199 -249
rect 199 -250 200 -249
rect 200 -250 201 -249
rect 201 -250 202 -249
rect 202 -250 203 -249
rect 203 -250 204 -249
rect 204 -250 205 -249
rect 205 -250 206 -249
rect 206 -250 207 -249
rect 207 -250 208 -249
rect 208 -250 209 -249
rect 209 -250 210 -249
rect 210 -250 211 -249
rect 211 -250 212 -249
rect 212 -250 213 -249
rect 213 -250 214 -249
rect 214 -250 215 -249
rect 215 -250 216 -249
rect 216 -250 217 -249
rect 217 -250 218 -249
rect 218 -250 219 -249
rect 219 -250 220 -249
rect 220 -250 221 -249
rect 221 -250 222 -249
rect 222 -250 223 -249
rect 223 -250 224 -249
rect 224 -250 225 -249
rect 225 -250 226 -249
rect 226 -250 227 -249
rect 227 -250 228 -249
rect 228 -250 229 -249
rect 229 -250 230 -249
rect 230 -250 231 -249
rect 231 -250 232 -249
rect 232 -250 233 -249
rect 233 -250 234 -249
rect 234 -250 235 -249
rect 235 -250 236 -249
rect 236 -250 237 -249
rect 237 -250 238 -249
rect 238 -250 239 -249
rect 239 -250 240 -249
rect 240 -250 241 -249
rect 241 -250 242 -249
rect 242 -250 243 -249
rect 243 -250 244 -249
rect 244 -250 245 -249
rect 245 -250 246 -249
rect 246 -250 247 -249
rect 247 -250 248 -249
rect 248 -250 249 -249
rect 249 -250 250 -249
rect 250 -250 251 -249
rect 251 -250 252 -249
rect 252 -250 253 -249
rect 253 -250 254 -249
rect 254 -250 255 -249
rect 255 -250 256 -249
rect 256 -250 257 -249
rect 257 -250 258 -249
rect 258 -250 259 -249
rect 259 -250 260 -249
rect 260 -250 261 -249
rect 261 -250 262 -249
rect 262 -250 263 -249
rect 263 -250 264 -249
rect 264 -250 265 -249
rect 265 -250 266 -249
rect 266 -250 267 -249
rect 267 -250 268 -249
rect 268 -250 269 -249
rect 269 -250 270 -249
rect 270 -250 271 -249
rect 271 -250 272 -249
rect 272 -250 273 -249
rect 273 -250 274 -249
rect 274 -250 275 -249
rect 275 -250 276 -249
rect 276 -250 277 -249
rect 277 -250 278 -249
rect 278 -250 279 -249
rect 279 -250 280 -249
rect 280 -250 281 -249
rect 281 -250 282 -249
rect 282 -250 283 -249
rect 283 -250 284 -249
rect 284 -250 285 -249
rect 285 -250 286 -249
rect 286 -250 287 -249
rect 287 -250 288 -249
rect 288 -250 289 -249
rect 289 -250 290 -249
rect 290 -250 291 -249
rect 291 -250 292 -249
rect 292 -250 293 -249
rect 293 -250 294 -249
rect 294 -250 295 -249
rect 295 -250 296 -249
rect 296 -250 297 -249
rect 297 -250 298 -249
rect 298 -250 299 -249
rect 299 -250 300 -249
rect 300 -250 301 -249
rect 301 -250 302 -249
rect 302 -250 303 -249
rect 303 -250 304 -249
rect 304 -250 305 -249
rect 305 -250 306 -249
rect 306 -250 307 -249
rect 307 -250 308 -249
rect 308 -250 309 -249
rect 309 -250 310 -249
rect 310 -250 311 -249
rect 311 -250 312 -249
rect 312 -250 313 -249
rect 313 -250 314 -249
rect 314 -250 315 -249
rect 315 -250 316 -249
rect 316 -250 317 -249
rect 317 -250 318 -249
rect 318 -250 319 -249
rect 319 -250 320 -249
rect 320 -250 321 -249
rect 321 -250 322 -249
rect 322 -250 323 -249
rect 323 -250 324 -249
rect 324 -250 325 -249
rect 325 -250 326 -249
rect 326 -250 327 -249
rect 327 -250 328 -249
rect 328 -250 329 -249
rect 329 -250 330 -249
rect 330 -250 331 -249
rect 331 -250 332 -249
rect 332 -250 333 -249
rect 333 -250 334 -249
rect 334 -250 335 -249
rect 335 -250 336 -249
rect 336 -250 337 -249
rect 337 -250 338 -249
rect 338 -250 339 -249
rect 339 -250 340 -249
rect 340 -250 341 -249
rect 341 -250 342 -249
rect 342 -250 343 -249
rect 343 -250 344 -249
rect 344 -250 345 -249
rect 345 -250 346 -249
rect 346 -250 347 -249
rect 347 -250 348 -249
rect 348 -250 349 -249
rect 349 -250 350 -249
rect 350 -250 351 -249
rect 351 -250 352 -249
rect 352 -250 353 -249
rect 353 -250 354 -249
rect 354 -250 355 -249
rect 355 -250 356 -249
rect 356 -250 357 -249
rect 357 -250 358 -249
rect 358 -250 359 -249
rect 359 -250 360 -249
rect 360 -250 361 -249
rect 361 -250 362 -249
rect 362 -250 363 -249
rect 363 -250 364 -249
rect 364 -250 365 -249
rect 365 -250 366 -249
rect 366 -250 367 -249
rect 367 -250 368 -249
rect 368 -250 369 -249
rect 369 -250 370 -249
rect 370 -250 371 -249
rect 371 -250 372 -249
rect 372 -250 373 -249
rect 373 -250 374 -249
rect 374 -250 375 -249
rect 375 -250 376 -249
rect 376 -250 377 -249
rect 377 -250 378 -249
rect 378 -250 379 -249
rect 379 -250 380 -249
rect 380 -250 381 -249
rect 381 -250 382 -249
rect 382 -250 383 -249
rect 383 -250 384 -249
rect 384 -250 385 -249
rect 385 -250 386 -249
rect 386 -250 387 -249
rect 387 -250 388 -249
rect 388 -250 389 -249
rect 389 -250 390 -249
rect 390 -250 391 -249
rect 391 -250 392 -249
rect 392 -250 393 -249
rect 393 -250 394 -249
rect 394 -250 395 -249
rect 395 -250 396 -249
rect 396 -250 397 -249
rect 397 -250 398 -249
rect 398 -250 399 -249
rect 399 -250 400 -249
rect 400 -250 401 -249
rect 401 -250 402 -249
rect 402 -250 403 -249
rect 403 -250 404 -249
rect 404 -250 405 -249
rect 405 -250 406 -249
rect 406 -250 407 -249
rect 407 -250 408 -249
rect 408 -250 409 -249
rect 409 -250 410 -249
rect 410 -250 411 -249
rect 411 -250 412 -249
rect 412 -250 413 -249
rect 413 -250 414 -249
rect 414 -250 415 -249
rect 415 -250 416 -249
rect 416 -250 417 -249
rect 417 -250 418 -249
rect 418 -250 419 -249
rect 419 -250 420 -249
rect 420 -250 421 -249
rect 421 -250 422 -249
rect 422 -250 423 -249
rect 423 -250 424 -249
rect 424 -250 425 -249
rect 425 -250 426 -249
rect 426 -250 427 -249
rect 427 -250 428 -249
rect 428 -250 429 -249
rect 429 -250 430 -249
rect 430 -250 431 -249
rect 431 -250 432 -249
rect 432 -250 433 -249
rect 433 -250 434 -249
rect 434 -250 435 -249
rect 435 -250 436 -249
rect 436 -250 437 -249
rect 437 -250 438 -249
rect 438 -250 439 -249
rect 439 -250 440 -249
rect 440 -250 441 -249
rect 441 -250 442 -249
rect 442 -250 443 -249
rect 443 -250 444 -249
rect 444 -250 445 -249
rect 445 -250 446 -249
rect 446 -250 447 -249
rect 447 -250 448 -249
rect 448 -250 449 -249
rect 449 -250 450 -249
rect 450 -250 451 -249
rect 451 -250 452 -249
rect 452 -250 453 -249
rect 453 -250 454 -249
rect 454 -250 455 -249
rect 455 -250 456 -249
rect 456 -250 457 -249
rect 457 -250 458 -249
rect 458 -250 459 -249
rect 459 -250 460 -249
rect 460 -250 461 -249
rect 461 -250 462 -249
rect 462 -250 463 -249
rect 463 -250 464 -249
rect 464 -250 465 -249
rect 465 -250 466 -249
rect 466 -250 467 -249
rect 467 -250 468 -249
rect 468 -250 469 -249
rect 469 -250 470 -249
rect 470 -250 471 -249
rect 471 -250 472 -249
rect 472 -250 473 -249
rect 473 -250 474 -249
rect 474 -250 475 -249
rect 475 -250 476 -249
rect 476 -250 477 -249
rect 477 -250 478 -249
rect 478 -250 479 -249
rect 479 -250 480 -249
rect 2 -251 3 -250
rect 3 -251 4 -250
rect 4 -251 5 -250
rect 5 -251 6 -250
rect 6 -251 7 -250
rect 7 -251 8 -250
rect 8 -251 9 -250
rect 9 -251 10 -250
rect 10 -251 11 -250
rect 11 -251 12 -250
rect 12 -251 13 -250
rect 13 -251 14 -250
rect 14 -251 15 -250
rect 15 -251 16 -250
rect 16 -251 17 -250
rect 17 -251 18 -250
rect 18 -251 19 -250
rect 19 -251 20 -250
rect 20 -251 21 -250
rect 21 -251 22 -250
rect 22 -251 23 -250
rect 23 -251 24 -250
rect 24 -251 25 -250
rect 25 -251 26 -250
rect 26 -251 27 -250
rect 27 -251 28 -250
rect 28 -251 29 -250
rect 29 -251 30 -250
rect 30 -251 31 -250
rect 31 -251 32 -250
rect 32 -251 33 -250
rect 33 -251 34 -250
rect 34 -251 35 -250
rect 35 -251 36 -250
rect 36 -251 37 -250
rect 37 -251 38 -250
rect 38 -251 39 -250
rect 39 -251 40 -250
rect 40 -251 41 -250
rect 41 -251 42 -250
rect 42 -251 43 -250
rect 43 -251 44 -250
rect 44 -251 45 -250
rect 45 -251 46 -250
rect 46 -251 47 -250
rect 47 -251 48 -250
rect 48 -251 49 -250
rect 49 -251 50 -250
rect 50 -251 51 -250
rect 51 -251 52 -250
rect 52 -251 53 -250
rect 53 -251 54 -250
rect 54 -251 55 -250
rect 55 -251 56 -250
rect 56 -251 57 -250
rect 57 -251 58 -250
rect 58 -251 59 -250
rect 59 -251 60 -250
rect 60 -251 61 -250
rect 61 -251 62 -250
rect 62 -251 63 -250
rect 63 -251 64 -250
rect 64 -251 65 -250
rect 65 -251 66 -250
rect 66 -251 67 -250
rect 67 -251 68 -250
rect 68 -251 69 -250
rect 69 -251 70 -250
rect 70 -251 71 -250
rect 71 -251 72 -250
rect 72 -251 73 -250
rect 73 -251 74 -250
rect 74 -251 75 -250
rect 75 -251 76 -250
rect 76 -251 77 -250
rect 77 -251 78 -250
rect 78 -251 79 -250
rect 79 -251 80 -250
rect 80 -251 81 -250
rect 81 -251 82 -250
rect 82 -251 83 -250
rect 83 -251 84 -250
rect 84 -251 85 -250
rect 85 -251 86 -250
rect 86 -251 87 -250
rect 87 -251 88 -250
rect 88 -251 89 -250
rect 89 -251 90 -250
rect 90 -251 91 -250
rect 91 -251 92 -250
rect 92 -251 93 -250
rect 93 -251 94 -250
rect 94 -251 95 -250
rect 95 -251 96 -250
rect 96 -251 97 -250
rect 97 -251 98 -250
rect 98 -251 99 -250
rect 99 -251 100 -250
rect 100 -251 101 -250
rect 101 -251 102 -250
rect 102 -251 103 -250
rect 103 -251 104 -250
rect 104 -251 105 -250
rect 105 -251 106 -250
rect 106 -251 107 -250
rect 107 -251 108 -250
rect 108 -251 109 -250
rect 109 -251 110 -250
rect 110 -251 111 -250
rect 111 -251 112 -250
rect 112 -251 113 -250
rect 113 -251 114 -250
rect 114 -251 115 -250
rect 115 -251 116 -250
rect 116 -251 117 -250
rect 117 -251 118 -250
rect 118 -251 119 -250
rect 119 -251 120 -250
rect 120 -251 121 -250
rect 121 -251 122 -250
rect 122 -251 123 -250
rect 123 -251 124 -250
rect 124 -251 125 -250
rect 125 -251 126 -250
rect 126 -251 127 -250
rect 127 -251 128 -250
rect 128 -251 129 -250
rect 129 -251 130 -250
rect 130 -251 131 -250
rect 131 -251 132 -250
rect 132 -251 133 -250
rect 133 -251 134 -250
rect 134 -251 135 -250
rect 135 -251 136 -250
rect 136 -251 137 -250
rect 137 -251 138 -250
rect 138 -251 139 -250
rect 139 -251 140 -250
rect 140 -251 141 -250
rect 141 -251 142 -250
rect 142 -251 143 -250
rect 143 -251 144 -250
rect 144 -251 145 -250
rect 145 -251 146 -250
rect 146 -251 147 -250
rect 147 -251 148 -250
rect 148 -251 149 -250
rect 149 -251 150 -250
rect 150 -251 151 -250
rect 151 -251 152 -250
rect 152 -251 153 -250
rect 153 -251 154 -250
rect 154 -251 155 -250
rect 155 -251 156 -250
rect 156 -251 157 -250
rect 157 -251 158 -250
rect 158 -251 159 -250
rect 159 -251 160 -250
rect 160 -251 161 -250
rect 161 -251 162 -250
rect 162 -251 163 -250
rect 163 -251 164 -250
rect 164 -251 165 -250
rect 165 -251 166 -250
rect 166 -251 167 -250
rect 167 -251 168 -250
rect 168 -251 169 -250
rect 169 -251 170 -250
rect 170 -251 171 -250
rect 171 -251 172 -250
rect 172 -251 173 -250
rect 173 -251 174 -250
rect 174 -251 175 -250
rect 175 -251 176 -250
rect 176 -251 177 -250
rect 177 -251 178 -250
rect 178 -251 179 -250
rect 179 -251 180 -250
rect 180 -251 181 -250
rect 181 -251 182 -250
rect 182 -251 183 -250
rect 183 -251 184 -250
rect 184 -251 185 -250
rect 185 -251 186 -250
rect 186 -251 187 -250
rect 187 -251 188 -250
rect 188 -251 189 -250
rect 189 -251 190 -250
rect 190 -251 191 -250
rect 191 -251 192 -250
rect 192 -251 193 -250
rect 193 -251 194 -250
rect 194 -251 195 -250
rect 195 -251 196 -250
rect 196 -251 197 -250
rect 197 -251 198 -250
rect 198 -251 199 -250
rect 199 -251 200 -250
rect 200 -251 201 -250
rect 201 -251 202 -250
rect 202 -251 203 -250
rect 203 -251 204 -250
rect 204 -251 205 -250
rect 205 -251 206 -250
rect 206 -251 207 -250
rect 207 -251 208 -250
rect 208 -251 209 -250
rect 209 -251 210 -250
rect 210 -251 211 -250
rect 211 -251 212 -250
rect 212 -251 213 -250
rect 213 -251 214 -250
rect 214 -251 215 -250
rect 215 -251 216 -250
rect 216 -251 217 -250
rect 217 -251 218 -250
rect 218 -251 219 -250
rect 219 -251 220 -250
rect 220 -251 221 -250
rect 221 -251 222 -250
rect 222 -251 223 -250
rect 223 -251 224 -250
rect 224 -251 225 -250
rect 225 -251 226 -250
rect 226 -251 227 -250
rect 227 -251 228 -250
rect 228 -251 229 -250
rect 229 -251 230 -250
rect 230 -251 231 -250
rect 231 -251 232 -250
rect 232 -251 233 -250
rect 233 -251 234 -250
rect 234 -251 235 -250
rect 235 -251 236 -250
rect 236 -251 237 -250
rect 237 -251 238 -250
rect 238 -251 239 -250
rect 239 -251 240 -250
rect 240 -251 241 -250
rect 241 -251 242 -250
rect 242 -251 243 -250
rect 243 -251 244 -250
rect 244 -251 245 -250
rect 245 -251 246 -250
rect 246 -251 247 -250
rect 247 -251 248 -250
rect 248 -251 249 -250
rect 249 -251 250 -250
rect 250 -251 251 -250
rect 251 -251 252 -250
rect 252 -251 253 -250
rect 253 -251 254 -250
rect 254 -251 255 -250
rect 255 -251 256 -250
rect 256 -251 257 -250
rect 257 -251 258 -250
rect 258 -251 259 -250
rect 259 -251 260 -250
rect 260 -251 261 -250
rect 261 -251 262 -250
rect 262 -251 263 -250
rect 263 -251 264 -250
rect 264 -251 265 -250
rect 265 -251 266 -250
rect 266 -251 267 -250
rect 267 -251 268 -250
rect 268 -251 269 -250
rect 269 -251 270 -250
rect 270 -251 271 -250
rect 271 -251 272 -250
rect 272 -251 273 -250
rect 273 -251 274 -250
rect 274 -251 275 -250
rect 275 -251 276 -250
rect 276 -251 277 -250
rect 277 -251 278 -250
rect 278 -251 279 -250
rect 279 -251 280 -250
rect 280 -251 281 -250
rect 281 -251 282 -250
rect 282 -251 283 -250
rect 283 -251 284 -250
rect 284 -251 285 -250
rect 285 -251 286 -250
rect 286 -251 287 -250
rect 287 -251 288 -250
rect 288 -251 289 -250
rect 289 -251 290 -250
rect 290 -251 291 -250
rect 291 -251 292 -250
rect 292 -251 293 -250
rect 293 -251 294 -250
rect 294 -251 295 -250
rect 295 -251 296 -250
rect 296 -251 297 -250
rect 297 -251 298 -250
rect 298 -251 299 -250
rect 299 -251 300 -250
rect 300 -251 301 -250
rect 301 -251 302 -250
rect 302 -251 303 -250
rect 303 -251 304 -250
rect 304 -251 305 -250
rect 305 -251 306 -250
rect 306 -251 307 -250
rect 307 -251 308 -250
rect 308 -251 309 -250
rect 309 -251 310 -250
rect 310 -251 311 -250
rect 311 -251 312 -250
rect 312 -251 313 -250
rect 313 -251 314 -250
rect 314 -251 315 -250
rect 315 -251 316 -250
rect 316 -251 317 -250
rect 317 -251 318 -250
rect 318 -251 319 -250
rect 319 -251 320 -250
rect 320 -251 321 -250
rect 321 -251 322 -250
rect 322 -251 323 -250
rect 323 -251 324 -250
rect 324 -251 325 -250
rect 325 -251 326 -250
rect 326 -251 327 -250
rect 327 -251 328 -250
rect 328 -251 329 -250
rect 329 -251 330 -250
rect 330 -251 331 -250
rect 331 -251 332 -250
rect 332 -251 333 -250
rect 333 -251 334 -250
rect 334 -251 335 -250
rect 335 -251 336 -250
rect 336 -251 337 -250
rect 337 -251 338 -250
rect 338 -251 339 -250
rect 339 -251 340 -250
rect 340 -251 341 -250
rect 341 -251 342 -250
rect 342 -251 343 -250
rect 343 -251 344 -250
rect 344 -251 345 -250
rect 345 -251 346 -250
rect 346 -251 347 -250
rect 347 -251 348 -250
rect 348 -251 349 -250
rect 349 -251 350 -250
rect 350 -251 351 -250
rect 351 -251 352 -250
rect 352 -251 353 -250
rect 353 -251 354 -250
rect 354 -251 355 -250
rect 355 -251 356 -250
rect 356 -251 357 -250
rect 357 -251 358 -250
rect 358 -251 359 -250
rect 359 -251 360 -250
rect 360 -251 361 -250
rect 361 -251 362 -250
rect 362 -251 363 -250
rect 363 -251 364 -250
rect 364 -251 365 -250
rect 365 -251 366 -250
rect 366 -251 367 -250
rect 367 -251 368 -250
rect 368 -251 369 -250
rect 369 -251 370 -250
rect 370 -251 371 -250
rect 371 -251 372 -250
rect 372 -251 373 -250
rect 373 -251 374 -250
rect 374 -251 375 -250
rect 375 -251 376 -250
rect 376 -251 377 -250
rect 377 -251 378 -250
rect 378 -251 379 -250
rect 379 -251 380 -250
rect 380 -251 381 -250
rect 381 -251 382 -250
rect 382 -251 383 -250
rect 383 -251 384 -250
rect 384 -251 385 -250
rect 385 -251 386 -250
rect 386 -251 387 -250
rect 387 -251 388 -250
rect 388 -251 389 -250
rect 389 -251 390 -250
rect 390 -251 391 -250
rect 391 -251 392 -250
rect 392 -251 393 -250
rect 393 -251 394 -250
rect 394 -251 395 -250
rect 395 -251 396 -250
rect 396 -251 397 -250
rect 397 -251 398 -250
rect 398 -251 399 -250
rect 399 -251 400 -250
rect 400 -251 401 -250
rect 401 -251 402 -250
rect 402 -251 403 -250
rect 403 -251 404 -250
rect 404 -251 405 -250
rect 405 -251 406 -250
rect 406 -251 407 -250
rect 407 -251 408 -250
rect 408 -251 409 -250
rect 409 -251 410 -250
rect 410 -251 411 -250
rect 411 -251 412 -250
rect 412 -251 413 -250
rect 413 -251 414 -250
rect 414 -251 415 -250
rect 415 -251 416 -250
rect 416 -251 417 -250
rect 417 -251 418 -250
rect 418 -251 419 -250
rect 419 -251 420 -250
rect 420 -251 421 -250
rect 421 -251 422 -250
rect 422 -251 423 -250
rect 423 -251 424 -250
rect 424 -251 425 -250
rect 425 -251 426 -250
rect 426 -251 427 -250
rect 427 -251 428 -250
rect 428 -251 429 -250
rect 429 -251 430 -250
rect 430 -251 431 -250
rect 431 -251 432 -250
rect 432 -251 433 -250
rect 433 -251 434 -250
rect 434 -251 435 -250
rect 435 -251 436 -250
rect 436 -251 437 -250
rect 437 -251 438 -250
rect 438 -251 439 -250
rect 439 -251 440 -250
rect 440 -251 441 -250
rect 441 -251 442 -250
rect 442 -251 443 -250
rect 443 -251 444 -250
rect 444 -251 445 -250
rect 445 -251 446 -250
rect 446 -251 447 -250
rect 447 -251 448 -250
rect 448 -251 449 -250
rect 449 -251 450 -250
rect 450 -251 451 -250
rect 451 -251 452 -250
rect 452 -251 453 -250
rect 453 -251 454 -250
rect 454 -251 455 -250
rect 455 -251 456 -250
rect 456 -251 457 -250
rect 457 -251 458 -250
rect 458 -251 459 -250
rect 459 -251 460 -250
rect 460 -251 461 -250
rect 461 -251 462 -250
rect 462 -251 463 -250
rect 463 -251 464 -250
rect 464 -251 465 -250
rect 465 -251 466 -250
rect 466 -251 467 -250
rect 467 -251 468 -250
rect 468 -251 469 -250
rect 469 -251 470 -250
rect 470 -251 471 -250
rect 471 -251 472 -250
rect 472 -251 473 -250
rect 473 -251 474 -250
rect 474 -251 475 -250
rect 475 -251 476 -250
rect 476 -251 477 -250
rect 477 -251 478 -250
rect 478 -251 479 -250
rect 479 -251 480 -250
rect 2 -252 3 -251
rect 3 -252 4 -251
rect 4 -252 5 -251
rect 5 -252 6 -251
rect 6 -252 7 -251
rect 7 -252 8 -251
rect 8 -252 9 -251
rect 9 -252 10 -251
rect 10 -252 11 -251
rect 11 -252 12 -251
rect 12 -252 13 -251
rect 13 -252 14 -251
rect 14 -252 15 -251
rect 15 -252 16 -251
rect 16 -252 17 -251
rect 17 -252 18 -251
rect 18 -252 19 -251
rect 19 -252 20 -251
rect 20 -252 21 -251
rect 21 -252 22 -251
rect 22 -252 23 -251
rect 23 -252 24 -251
rect 24 -252 25 -251
rect 25 -252 26 -251
rect 26 -252 27 -251
rect 27 -252 28 -251
rect 28 -252 29 -251
rect 29 -252 30 -251
rect 30 -252 31 -251
rect 31 -252 32 -251
rect 32 -252 33 -251
rect 33 -252 34 -251
rect 34 -252 35 -251
rect 35 -252 36 -251
rect 36 -252 37 -251
rect 37 -252 38 -251
rect 38 -252 39 -251
rect 39 -252 40 -251
rect 40 -252 41 -251
rect 41 -252 42 -251
rect 42 -252 43 -251
rect 43 -252 44 -251
rect 44 -252 45 -251
rect 45 -252 46 -251
rect 46 -252 47 -251
rect 47 -252 48 -251
rect 48 -252 49 -251
rect 49 -252 50 -251
rect 50 -252 51 -251
rect 51 -252 52 -251
rect 52 -252 53 -251
rect 53 -252 54 -251
rect 54 -252 55 -251
rect 55 -252 56 -251
rect 56 -252 57 -251
rect 57 -252 58 -251
rect 58 -252 59 -251
rect 59 -252 60 -251
rect 60 -252 61 -251
rect 61 -252 62 -251
rect 62 -252 63 -251
rect 63 -252 64 -251
rect 64 -252 65 -251
rect 65 -252 66 -251
rect 66 -252 67 -251
rect 67 -252 68 -251
rect 68 -252 69 -251
rect 69 -252 70 -251
rect 70 -252 71 -251
rect 71 -252 72 -251
rect 72 -252 73 -251
rect 73 -252 74 -251
rect 74 -252 75 -251
rect 75 -252 76 -251
rect 76 -252 77 -251
rect 77 -252 78 -251
rect 78 -252 79 -251
rect 79 -252 80 -251
rect 80 -252 81 -251
rect 81 -252 82 -251
rect 82 -252 83 -251
rect 83 -252 84 -251
rect 84 -252 85 -251
rect 85 -252 86 -251
rect 86 -252 87 -251
rect 87 -252 88 -251
rect 88 -252 89 -251
rect 89 -252 90 -251
rect 90 -252 91 -251
rect 91 -252 92 -251
rect 92 -252 93 -251
rect 93 -252 94 -251
rect 94 -252 95 -251
rect 95 -252 96 -251
rect 96 -252 97 -251
rect 97 -252 98 -251
rect 98 -252 99 -251
rect 99 -252 100 -251
rect 100 -252 101 -251
rect 101 -252 102 -251
rect 102 -252 103 -251
rect 103 -252 104 -251
rect 104 -252 105 -251
rect 105 -252 106 -251
rect 106 -252 107 -251
rect 107 -252 108 -251
rect 108 -252 109 -251
rect 109 -252 110 -251
rect 110 -252 111 -251
rect 111 -252 112 -251
rect 112 -252 113 -251
rect 113 -252 114 -251
rect 114 -252 115 -251
rect 115 -252 116 -251
rect 116 -252 117 -251
rect 117 -252 118 -251
rect 118 -252 119 -251
rect 119 -252 120 -251
rect 120 -252 121 -251
rect 121 -252 122 -251
rect 122 -252 123 -251
rect 123 -252 124 -251
rect 124 -252 125 -251
rect 125 -252 126 -251
rect 126 -252 127 -251
rect 127 -252 128 -251
rect 128 -252 129 -251
rect 129 -252 130 -251
rect 130 -252 131 -251
rect 131 -252 132 -251
rect 132 -252 133 -251
rect 133 -252 134 -251
rect 134 -252 135 -251
rect 135 -252 136 -251
rect 136 -252 137 -251
rect 137 -252 138 -251
rect 138 -252 139 -251
rect 139 -252 140 -251
rect 140 -252 141 -251
rect 141 -252 142 -251
rect 142 -252 143 -251
rect 143 -252 144 -251
rect 144 -252 145 -251
rect 145 -252 146 -251
rect 146 -252 147 -251
rect 147 -252 148 -251
rect 148 -252 149 -251
rect 149 -252 150 -251
rect 150 -252 151 -251
rect 151 -252 152 -251
rect 152 -252 153 -251
rect 153 -252 154 -251
rect 154 -252 155 -251
rect 155 -252 156 -251
rect 156 -252 157 -251
rect 157 -252 158 -251
rect 158 -252 159 -251
rect 159 -252 160 -251
rect 160 -252 161 -251
rect 161 -252 162 -251
rect 162 -252 163 -251
rect 163 -252 164 -251
rect 164 -252 165 -251
rect 165 -252 166 -251
rect 166 -252 167 -251
rect 167 -252 168 -251
rect 168 -252 169 -251
rect 169 -252 170 -251
rect 170 -252 171 -251
rect 171 -252 172 -251
rect 172 -252 173 -251
rect 173 -252 174 -251
rect 174 -252 175 -251
rect 175 -252 176 -251
rect 176 -252 177 -251
rect 177 -252 178 -251
rect 178 -252 179 -251
rect 179 -252 180 -251
rect 180 -252 181 -251
rect 181 -252 182 -251
rect 182 -252 183 -251
rect 183 -252 184 -251
rect 184 -252 185 -251
rect 185 -252 186 -251
rect 186 -252 187 -251
rect 187 -252 188 -251
rect 188 -252 189 -251
rect 189 -252 190 -251
rect 190 -252 191 -251
rect 191 -252 192 -251
rect 192 -252 193 -251
rect 193 -252 194 -251
rect 194 -252 195 -251
rect 195 -252 196 -251
rect 196 -252 197 -251
rect 197 -252 198 -251
rect 198 -252 199 -251
rect 199 -252 200 -251
rect 200 -252 201 -251
rect 201 -252 202 -251
rect 202 -252 203 -251
rect 203 -252 204 -251
rect 204 -252 205 -251
rect 205 -252 206 -251
rect 206 -252 207 -251
rect 207 -252 208 -251
rect 208 -252 209 -251
rect 209 -252 210 -251
rect 210 -252 211 -251
rect 211 -252 212 -251
rect 212 -252 213 -251
rect 213 -252 214 -251
rect 214 -252 215 -251
rect 215 -252 216 -251
rect 216 -252 217 -251
rect 217 -252 218 -251
rect 218 -252 219 -251
rect 219 -252 220 -251
rect 220 -252 221 -251
rect 221 -252 222 -251
rect 222 -252 223 -251
rect 223 -252 224 -251
rect 224 -252 225 -251
rect 225 -252 226 -251
rect 226 -252 227 -251
rect 227 -252 228 -251
rect 228 -252 229 -251
rect 229 -252 230 -251
rect 230 -252 231 -251
rect 231 -252 232 -251
rect 232 -252 233 -251
rect 233 -252 234 -251
rect 234 -252 235 -251
rect 235 -252 236 -251
rect 236 -252 237 -251
rect 237 -252 238 -251
rect 238 -252 239 -251
rect 239 -252 240 -251
rect 240 -252 241 -251
rect 241 -252 242 -251
rect 242 -252 243 -251
rect 243 -252 244 -251
rect 244 -252 245 -251
rect 245 -252 246 -251
rect 246 -252 247 -251
rect 247 -252 248 -251
rect 248 -252 249 -251
rect 249 -252 250 -251
rect 250 -252 251 -251
rect 251 -252 252 -251
rect 252 -252 253 -251
rect 253 -252 254 -251
rect 254 -252 255 -251
rect 255 -252 256 -251
rect 256 -252 257 -251
rect 257 -252 258 -251
rect 258 -252 259 -251
rect 259 -252 260 -251
rect 260 -252 261 -251
rect 261 -252 262 -251
rect 262 -252 263 -251
rect 263 -252 264 -251
rect 264 -252 265 -251
rect 265 -252 266 -251
rect 266 -252 267 -251
rect 267 -252 268 -251
rect 268 -252 269 -251
rect 269 -252 270 -251
rect 270 -252 271 -251
rect 271 -252 272 -251
rect 272 -252 273 -251
rect 273 -252 274 -251
rect 274 -252 275 -251
rect 275 -252 276 -251
rect 276 -252 277 -251
rect 277 -252 278 -251
rect 278 -252 279 -251
rect 279 -252 280 -251
rect 280 -252 281 -251
rect 281 -252 282 -251
rect 282 -252 283 -251
rect 283 -252 284 -251
rect 284 -252 285 -251
rect 285 -252 286 -251
rect 286 -252 287 -251
rect 287 -252 288 -251
rect 288 -252 289 -251
rect 289 -252 290 -251
rect 290 -252 291 -251
rect 291 -252 292 -251
rect 292 -252 293 -251
rect 293 -252 294 -251
rect 294 -252 295 -251
rect 295 -252 296 -251
rect 296 -252 297 -251
rect 297 -252 298 -251
rect 298 -252 299 -251
rect 299 -252 300 -251
rect 300 -252 301 -251
rect 301 -252 302 -251
rect 302 -252 303 -251
rect 303 -252 304 -251
rect 304 -252 305 -251
rect 305 -252 306 -251
rect 306 -252 307 -251
rect 307 -252 308 -251
rect 308 -252 309 -251
rect 309 -252 310 -251
rect 310 -252 311 -251
rect 311 -252 312 -251
rect 312 -252 313 -251
rect 313 -252 314 -251
rect 314 -252 315 -251
rect 315 -252 316 -251
rect 316 -252 317 -251
rect 317 -252 318 -251
rect 318 -252 319 -251
rect 319 -252 320 -251
rect 320 -252 321 -251
rect 321 -252 322 -251
rect 322 -252 323 -251
rect 323 -252 324 -251
rect 324 -252 325 -251
rect 325 -252 326 -251
rect 326 -252 327 -251
rect 327 -252 328 -251
rect 328 -252 329 -251
rect 329 -252 330 -251
rect 330 -252 331 -251
rect 331 -252 332 -251
rect 332 -252 333 -251
rect 333 -252 334 -251
rect 334 -252 335 -251
rect 335 -252 336 -251
rect 336 -252 337 -251
rect 337 -252 338 -251
rect 338 -252 339 -251
rect 339 -252 340 -251
rect 340 -252 341 -251
rect 341 -252 342 -251
rect 342 -252 343 -251
rect 343 -252 344 -251
rect 344 -252 345 -251
rect 345 -252 346 -251
rect 346 -252 347 -251
rect 347 -252 348 -251
rect 348 -252 349 -251
rect 349 -252 350 -251
rect 350 -252 351 -251
rect 351 -252 352 -251
rect 352 -252 353 -251
rect 353 -252 354 -251
rect 354 -252 355 -251
rect 355 -252 356 -251
rect 356 -252 357 -251
rect 357 -252 358 -251
rect 358 -252 359 -251
rect 359 -252 360 -251
rect 360 -252 361 -251
rect 361 -252 362 -251
rect 362 -252 363 -251
rect 363 -252 364 -251
rect 364 -252 365 -251
rect 365 -252 366 -251
rect 366 -252 367 -251
rect 367 -252 368 -251
rect 368 -252 369 -251
rect 369 -252 370 -251
rect 370 -252 371 -251
rect 371 -252 372 -251
rect 372 -252 373 -251
rect 373 -252 374 -251
rect 374 -252 375 -251
rect 375 -252 376 -251
rect 376 -252 377 -251
rect 377 -252 378 -251
rect 378 -252 379 -251
rect 379 -252 380 -251
rect 380 -252 381 -251
rect 381 -252 382 -251
rect 382 -252 383 -251
rect 383 -252 384 -251
rect 384 -252 385 -251
rect 385 -252 386 -251
rect 386 -252 387 -251
rect 387 -252 388 -251
rect 388 -252 389 -251
rect 389 -252 390 -251
rect 390 -252 391 -251
rect 391 -252 392 -251
rect 392 -252 393 -251
rect 393 -252 394 -251
rect 394 -252 395 -251
rect 395 -252 396 -251
rect 396 -252 397 -251
rect 397 -252 398 -251
rect 398 -252 399 -251
rect 399 -252 400 -251
rect 400 -252 401 -251
rect 401 -252 402 -251
rect 402 -252 403 -251
rect 403 -252 404 -251
rect 404 -252 405 -251
rect 405 -252 406 -251
rect 406 -252 407 -251
rect 407 -252 408 -251
rect 408 -252 409 -251
rect 409 -252 410 -251
rect 410 -252 411 -251
rect 411 -252 412 -251
rect 412 -252 413 -251
rect 413 -252 414 -251
rect 414 -252 415 -251
rect 415 -252 416 -251
rect 416 -252 417 -251
rect 417 -252 418 -251
rect 418 -252 419 -251
rect 419 -252 420 -251
rect 420 -252 421 -251
rect 421 -252 422 -251
rect 422 -252 423 -251
rect 423 -252 424 -251
rect 424 -252 425 -251
rect 425 -252 426 -251
rect 426 -252 427 -251
rect 427 -252 428 -251
rect 428 -252 429 -251
rect 429 -252 430 -251
rect 430 -252 431 -251
rect 431 -252 432 -251
rect 432 -252 433 -251
rect 433 -252 434 -251
rect 434 -252 435 -251
rect 435 -252 436 -251
rect 436 -252 437 -251
rect 437 -252 438 -251
rect 438 -252 439 -251
rect 439 -252 440 -251
rect 440 -252 441 -251
rect 441 -252 442 -251
rect 442 -252 443 -251
rect 443 -252 444 -251
rect 444 -252 445 -251
rect 445 -252 446 -251
rect 446 -252 447 -251
rect 447 -252 448 -251
rect 448 -252 449 -251
rect 449 -252 450 -251
rect 450 -252 451 -251
rect 451 -252 452 -251
rect 452 -252 453 -251
rect 453 -252 454 -251
rect 454 -252 455 -251
rect 455 -252 456 -251
rect 456 -252 457 -251
rect 457 -252 458 -251
rect 458 -252 459 -251
rect 459 -252 460 -251
rect 460 -252 461 -251
rect 461 -252 462 -251
rect 462 -252 463 -251
rect 463 -252 464 -251
rect 464 -252 465 -251
rect 465 -252 466 -251
rect 466 -252 467 -251
rect 467 -252 468 -251
rect 468 -252 469 -251
rect 469 -252 470 -251
rect 470 -252 471 -251
rect 471 -252 472 -251
rect 472 -252 473 -251
rect 473 -252 474 -251
rect 474 -252 475 -251
rect 475 -252 476 -251
rect 476 -252 477 -251
rect 477 -252 478 -251
rect 478 -252 479 -251
rect 479 -252 480 -251
<< end >>