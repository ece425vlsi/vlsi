magic
tech scmos
timestamp 1492531947
<< m2contact >>
rect 593 196 597 200
rect 30 167 34 171
rect 110 167 114 171
rect 190 167 194 171
rect 270 167 274 171
rect 350 167 354 171
rect 430 167 434 171
rect 510 167 514 171
rect 593 168 597 172
rect 593 140 597 144
rect 593 112 597 116
rect 593 84 597 88
rect 593 56 597 60
rect 198 42 202 46
rect 270 42 274 46
rect 593 28 597 32
rect 593 0 597 4
rect 619 0 623 4
rect 641 0 645 4
rect 663 0 667 4
rect 685 0 689 4
rect 707 0 711 4
rect 729 0 733 4
rect 751 0 755 4
<< metal2 >>
rect 550 200 555 201
rect 554 196 555 200
rect 70 108 74 163
rect 6 -59 10 46
rect 38 -50 42 46
rect 45 32 49 104
rect 150 78 154 163
rect 230 87 234 163
rect 310 96 314 163
rect 390 105 394 163
rect 470 159 474 179
rect 550 159 555 196
rect 579 172 583 179
rect 572 105 576 140
rect 581 92 585 112
rect 559 60 563 74
rect 70 -41 74 46
rect 102 -32 106 46
rect 134 -23 138 46
rect 166 -14 170 46
rect 198 -5 202 42
rect 280 4 284 42
rect 619 -5 623 0
rect 641 -14 645 0
rect 663 -23 667 0
rect 685 -32 689 0
rect 707 -41 711 0
rect 729 -50 733 0
rect 751 -59 755 0
<< m3contact >>
rect 550 196 554 200
rect 593 196 597 200
rect 470 179 474 183
rect 45 104 49 108
rect 70 104 74 108
rect 579 179 583 183
rect 579 168 583 172
rect 593 168 597 172
rect 390 101 394 105
rect 572 140 576 144
rect 593 140 597 144
rect 572 101 576 105
rect 581 112 585 116
rect 593 112 597 116
rect 310 92 314 96
rect 230 83 234 87
rect 593 84 597 88
rect 150 74 154 78
rect 559 74 563 78
rect 559 56 563 60
rect 593 56 597 60
rect 45 28 49 32
rect 270 42 274 46
rect 280 42 284 46
rect 593 28 597 32
rect 280 0 284 4
rect 593 0 597 4
rect 198 -9 202 -5
rect 619 -9 623 -5
rect 166 -18 170 -14
rect 641 -18 645 -14
rect 134 -27 138 -23
rect 663 -27 667 -23
rect 102 -36 106 -32
rect 685 -36 689 -32
rect 70 -45 74 -41
rect 707 -45 711 -41
rect 38 -54 42 -50
rect 729 -54 733 -50
rect 6 -63 10 -59
rect 751 -63 755 -59
<< metal3 >>
rect 549 200 598 201
rect 549 196 550 200
rect 554 196 593 200
rect 597 196 598 200
rect 549 195 598 196
rect 469 183 584 184
rect 469 179 470 183
rect 474 179 579 183
rect 583 179 584 183
rect 469 178 584 179
rect 578 172 598 173
rect 578 168 579 172
rect 583 168 593 172
rect 597 168 598 172
rect 578 167 598 168
rect 571 144 598 145
rect 571 140 572 144
rect 576 140 593 144
rect 597 140 598 144
rect 571 139 598 140
rect 580 116 598 117
rect 580 112 581 116
rect 585 112 593 116
rect 597 112 598 116
rect 580 111 598 112
rect 44 108 75 109
rect 44 104 45 108
rect 49 104 70 108
rect 74 104 75 108
rect 44 103 75 104
rect 389 105 577 106
rect 389 101 390 105
rect 394 101 572 105
rect 576 101 577 105
rect 389 100 577 101
rect 309 96 586 97
rect 309 92 310 96
rect 314 92 586 96
rect 309 91 586 92
rect 592 88 598 89
rect 229 87 593 88
rect 229 83 230 87
rect 234 84 593 87
rect 597 84 598 88
rect 234 83 598 84
rect 229 82 598 83
rect 149 78 564 79
rect 149 74 150 78
rect 154 74 559 78
rect 563 74 564 78
rect 149 73 564 74
rect 558 60 598 61
rect 558 56 559 60
rect 563 56 593 60
rect 597 56 598 60
rect 558 55 598 56
rect 269 46 285 47
rect 269 42 270 46
rect 274 42 280 46
rect 284 42 285 46
rect 269 41 285 42
rect 44 32 598 33
rect 44 28 45 32
rect 49 28 593 32
rect 597 28 598 32
rect 44 27 598 28
rect 279 4 598 5
rect 279 0 280 4
rect 284 0 593 4
rect 597 0 598 4
rect 279 -1 598 0
rect 197 -5 624 -4
rect 197 -9 198 -5
rect 202 -9 619 -5
rect 623 -9 624 -5
rect 197 -10 624 -9
rect 165 -14 646 -13
rect 165 -18 166 -14
rect 170 -18 641 -14
rect 645 -18 646 -14
rect 165 -19 646 -18
rect 133 -23 668 -22
rect 133 -27 134 -23
rect 138 -27 663 -23
rect 667 -27 668 -23
rect 133 -28 668 -27
rect 101 -32 690 -31
rect 101 -36 102 -32
rect 106 -36 685 -32
rect 689 -36 690 -32
rect 101 -37 690 -36
rect 69 -41 712 -40
rect 69 -45 70 -41
rect 74 -45 707 -41
rect 711 -45 712 -41
rect 69 -46 712 -45
rect 37 -50 734 -49
rect 37 -54 38 -50
rect 42 -54 729 -50
rect 733 -54 734 -50
rect 37 -55 734 -54
rect 5 -59 756 -58
rect 5 -63 6 -59
rect 10 -63 751 -59
rect 755 -63 756 -59
rect 5 -64 756 -63
use source_gen_7_0  source_gen_7_0_0
timestamp 1492528143
transform 1 0 0 0 1 0
box 0 0 773 224
<< end >>
