magic
tech scmos
timestamp 1488311656
<< m2contact >>
rect -7 -2 7 2
<< end >>
